module Mesh( // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177818.2]
  input         clock, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177819.4]
  input  [7:0]  io_in_a_0_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [7:0]  io_in_a_1_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [7:0]  io_in_a_2_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [7:0]  io_in_a_3_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [7:0]  io_in_a_4_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [7:0]  io_in_a_5_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [7:0]  io_in_a_6_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [7:0]  io_in_a_7_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [7:0]  io_in_d_0_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [7:0]  io_in_d_1_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [7:0]  io_in_d_2_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [7:0]  io_in_d_3_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [7:0]  io_in_d_4_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [7:0]  io_in_d_5_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [7:0]  io_in_d_6_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [7:0]  io_in_d_7_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [7:0]  io_in_b_0_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [7:0]  io_in_b_1_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [7:0]  io_in_b_2_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [7:0]  io_in_b_3_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [7:0]  io_in_b_4_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [7:0]  io_in_b_5_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [7:0]  io_in_b_6_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [7:0]  io_in_b_7_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input         io_in_control_0_0_propagate, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [5:0]  io_in_control_0_0_shift, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input         io_in_control_1_0_propagate, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [5:0]  io_in_control_1_0_shift, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input         io_in_control_2_0_propagate, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [5:0]  io_in_control_2_0_shift, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input         io_in_control_3_0_propagate, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [5:0]  io_in_control_3_0_shift, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input         io_in_control_4_0_propagate, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [5:0]  io_in_control_4_0_shift, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input         io_in_control_5_0_propagate, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [5:0]  io_in_control_5_0_shift, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input         io_in_control_6_0_propagate, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [5:0]  io_in_control_6_0_shift, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input         io_in_control_7_0_propagate, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input  [5:0]  io_in_control_7_0_shift, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  output reg [18:0] io_out_c_0_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  output reg [18:0] io_out_c_1_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  output reg [18:0] io_out_c_2_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  output reg [18:0] io_out_c_3_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  output reg [18:0] io_out_c_4_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  output reg [18:0] io_out_c_5_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  output reg [18:0] io_out_c_6_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  output reg [18:0] io_out_c_7_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  output [18:0] io_out_b_0_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  output [18:0] io_out_b_1_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  output [18:0] io_out_b_2_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  output [18:0] io_out_b_3_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  output [18:0] io_out_b_4_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  output [18:0] io_out_b_5_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  output [18:0] io_out_b_6_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  output [18:0] io_out_b_7_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input         io_in_valid_0_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input         io_in_valid_1_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input         io_in_valid_2_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input         io_in_valid_3_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input         io_in_valid_4_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input         io_in_valid_5_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input         io_in_valid_6_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  input         io_in_valid_7_0, // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
  output reg       io_out_valid_0_0 // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177821.4]
);


`include "parameters.v"

  wire  mesh_0_0_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177823.4]
  wire [7:0] mesh_0_0_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177823.4]
  wire [18:0] mesh_0_0_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177823.4]
  wire [18:0] mesh_0_0_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177823.4]
  wire  mesh_0_0_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177823.4]
  wire [5:0] mesh_0_0_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177823.4]
  wire [7:0] mesh_0_0_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177823.4]
  wire [(dbits-1):0] mesh_0_0_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177823.4]
  wire [18:0] mesh_0_0_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177823.4]
  wire  mesh_0_0_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177823.4]
  wire [5:0] mesh_0_0_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177823.4]
  wire  mesh_0_0_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177823.4]
  wire  mesh_0_0_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177823.4]
  wire  mesh_0_1_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177826.4]
  wire [7:0] mesh_0_1_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177826.4]
  wire [18:0] mesh_0_1_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177826.4]
  wire [18:0] mesh_0_1_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177826.4]
  wire  mesh_0_1_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177826.4]
  wire [5:0] mesh_0_1_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177826.4]
  wire [7:0] mesh_0_1_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177826.4]
  wire [(dbits-1):0] mesh_0_1_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177826.4]
  wire [18:0] mesh_0_1_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177826.4]
  wire  mesh_0_1_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177826.4]
  wire [5:0] mesh_0_1_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177826.4]
  wire  mesh_0_1_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177826.4]
  wire  mesh_0_1_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177826.4]
  wire  mesh_0_2_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177829.4]
  wire [7:0] mesh_0_2_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177829.4]
  wire [18:0] mesh_0_2_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177829.4]
  wire [18:0] mesh_0_2_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177829.4]
  wire  mesh_0_2_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177829.4]
  wire [5:0] mesh_0_2_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177829.4]
  wire [7:0] mesh_0_2_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177829.4]
  wire [(dbits-1):0] mesh_0_2_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177829.4]
  wire [18:0] mesh_0_2_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177829.4]
  wire  mesh_0_2_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177829.4]
  wire [5:0] mesh_0_2_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177829.4]
  wire  mesh_0_2_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177829.4]
  wire  mesh_0_2_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177829.4]
  wire  mesh_0_3_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177832.4]
  wire [7:0] mesh_0_3_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177832.4]
  wire [18:0] mesh_0_3_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177832.4]
  wire [18:0] mesh_0_3_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177832.4]
  wire  mesh_0_3_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177832.4]
  wire [5:0] mesh_0_3_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177832.4]
  wire [7:0] mesh_0_3_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177832.4]
  wire [(dbits-1):0] mesh_0_3_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177832.4]
  wire [18:0] mesh_0_3_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177832.4]
  wire  mesh_0_3_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177832.4]
  wire [5:0] mesh_0_3_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177832.4]
  wire  mesh_0_3_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177832.4]
  wire  mesh_0_3_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177832.4]
  wire  mesh_0_4_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177835.4]
  wire [7:0] mesh_0_4_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177835.4]
  wire [18:0] mesh_0_4_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177835.4]
  wire [18:0] mesh_0_4_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177835.4]
  wire  mesh_0_4_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177835.4]
  wire [5:0] mesh_0_4_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177835.4]
  wire [7:0] mesh_0_4_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177835.4]
  wire [(dbits-1):0] mesh_0_4_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177835.4]
  wire [18:0] mesh_0_4_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177835.4]
  wire  mesh_0_4_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177835.4]
  wire [5:0] mesh_0_4_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177835.4]
  wire  mesh_0_4_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177835.4]
  wire  mesh_0_4_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177835.4]
  wire  mesh_0_5_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177838.4]
  wire [7:0] mesh_0_5_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177838.4]
  wire [18:0] mesh_0_5_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177838.4]
  wire [18:0] mesh_0_5_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177838.4]
  wire  mesh_0_5_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177838.4]
  wire [5:0] mesh_0_5_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177838.4]
  wire [7:0] mesh_0_5_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177838.4]
  wire [(dbits-1):0] mesh_0_5_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177838.4]
  wire [18:0] mesh_0_5_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177838.4]
  wire  mesh_0_5_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177838.4]
  wire [5:0] mesh_0_5_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177838.4]
  wire  mesh_0_5_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177838.4]
  wire  mesh_0_5_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177838.4]
  wire  mesh_0_6_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177841.4]
  wire [7:0] mesh_0_6_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177841.4]
  wire [18:0] mesh_0_6_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177841.4]
  wire [18:0] mesh_0_6_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177841.4]
  wire  mesh_0_6_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177841.4]
  wire [5:0] mesh_0_6_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177841.4]
  wire [7:0] mesh_0_6_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177841.4]
  wire [(dbits-1):0] mesh_0_6_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177841.4]
  wire [18:0] mesh_0_6_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177841.4]
  wire  mesh_0_6_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177841.4]
  wire [5:0] mesh_0_6_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177841.4]
  wire  mesh_0_6_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177841.4]
  wire  mesh_0_6_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177841.4]
  wire  mesh_0_7_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177844.4]
  wire [7:0] mesh_0_7_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177844.4]
  wire [18:0] mesh_0_7_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177844.4]
  wire [18:0] mesh_0_7_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177844.4]
  wire  mesh_0_7_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177844.4]
  wire [5:0] mesh_0_7_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177844.4]
  wire [7:0] mesh_0_7_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177844.4]
  wire [(dbits-1):0] mesh_0_7_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177844.4]
  wire [18:0] mesh_0_7_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177844.4]
  wire  mesh_0_7_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177844.4]
  wire [5:0] mesh_0_7_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177844.4]
  wire  mesh_0_7_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177844.4]
  wire  mesh_0_7_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177844.4]
  wire  mesh_1_0_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177847.4]
  wire [7:0] mesh_1_0_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177847.4]
  wire [18:0] mesh_1_0_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177847.4]
  wire [(dbits-1):0] mesh_1_0_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177847.4]
  wire  mesh_1_0_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177847.4]
  wire [5:0] mesh_1_0_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177847.4]
  wire [7:0] mesh_1_0_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177847.4]
  wire [(dbits-1):0] mesh_1_0_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177847.4]
  wire [18:0] mesh_1_0_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177847.4]
  wire  mesh_1_0_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177847.4]
  wire [5:0] mesh_1_0_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177847.4]
  wire  mesh_1_0_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177847.4]
  wire  mesh_1_0_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177847.4]
  wire  mesh_1_1_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177850.4]
  wire [7:0] mesh_1_1_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177850.4]
  wire [18:0] mesh_1_1_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177850.4]
  wire [(dbits-1):0] mesh_1_1_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177850.4]
  wire  mesh_1_1_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177850.4]
  wire [5:0] mesh_1_1_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177850.4]
  wire [7:0] mesh_1_1_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177850.4]
  wire [(dbits-1):0] mesh_1_1_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177850.4]
  wire [18:0] mesh_1_1_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177850.4]
  wire  mesh_1_1_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177850.4]
  wire [5:0] mesh_1_1_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177850.4]
  wire  mesh_1_1_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177850.4]
  wire  mesh_1_1_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177850.4]
  wire  mesh_1_2_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177853.4]
  wire [7:0] mesh_1_2_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177853.4]
  wire [18:0] mesh_1_2_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177853.4]
  wire [(dbits-1):0] mesh_1_2_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177853.4]
  wire  mesh_1_2_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177853.4]
  wire [5:0] mesh_1_2_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177853.4]
  wire [7:0] mesh_1_2_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177853.4]
  wire [(dbits-1):0] mesh_1_2_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177853.4]
  wire [18:0] mesh_1_2_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177853.4]
  wire  mesh_1_2_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177853.4]
  wire [5:0] mesh_1_2_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177853.4]
  wire  mesh_1_2_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177853.4]
  wire  mesh_1_2_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177853.4]
  wire  mesh_1_3_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177856.4]
  wire [7:0] mesh_1_3_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177856.4]
  wire [18:0] mesh_1_3_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177856.4]
  wire [(dbits-1):0] mesh_1_3_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177856.4]
  wire  mesh_1_3_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177856.4]
  wire [5:0] mesh_1_3_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177856.4]
  wire [7:0] mesh_1_3_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177856.4]
  wire [(dbits-1):0] mesh_1_3_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177856.4]
  wire [18:0] mesh_1_3_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177856.4]
  wire  mesh_1_3_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177856.4]
  wire [5:0] mesh_1_3_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177856.4]
  wire  mesh_1_3_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177856.4]
  wire  mesh_1_3_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177856.4]
  wire  mesh_1_4_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177859.4]
  wire [7:0] mesh_1_4_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177859.4]
  wire [18:0] mesh_1_4_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177859.4]
  wire [(dbits-1):0] mesh_1_4_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177859.4]
  wire  mesh_1_4_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177859.4]
  wire [5:0] mesh_1_4_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177859.4]
  wire [7:0] mesh_1_4_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177859.4]
  wire [(dbits-1):0] mesh_1_4_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177859.4]
  wire [18:0] mesh_1_4_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177859.4]
  wire  mesh_1_4_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177859.4]
  wire [5:0] mesh_1_4_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177859.4]
  wire  mesh_1_4_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177859.4]
  wire  mesh_1_4_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177859.4]
  wire  mesh_1_5_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177862.4]
  wire [7:0] mesh_1_5_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177862.4]
  wire [18:0] mesh_1_5_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177862.4]
  wire [(dbits-1):0] mesh_1_5_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177862.4]
  wire  mesh_1_5_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177862.4]
  wire [5:0] mesh_1_5_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177862.4]
  wire [7:0] mesh_1_5_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177862.4]
  wire [(dbits-1):0] mesh_1_5_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177862.4]
  wire [18:0] mesh_1_5_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177862.4]
  wire  mesh_1_5_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177862.4]
  wire [5:0] mesh_1_5_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177862.4]
  wire  mesh_1_5_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177862.4]
  wire  mesh_1_5_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177862.4]
  wire  mesh_1_6_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177865.4]
  wire [7:0] mesh_1_6_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177865.4]
  wire [18:0] mesh_1_6_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177865.4]
  wire [(dbits-1):0] mesh_1_6_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177865.4]
  wire  mesh_1_6_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177865.4]
  wire [5:0] mesh_1_6_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177865.4]
  wire [7:0] mesh_1_6_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177865.4]
  wire [(dbits-1):0] mesh_1_6_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177865.4]
  wire [18:0] mesh_1_6_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177865.4]
  wire  mesh_1_6_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177865.4]
  wire [5:0] mesh_1_6_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177865.4]
  wire  mesh_1_6_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177865.4]
  wire  mesh_1_6_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177865.4]
  wire  mesh_1_7_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177868.4]
  wire [7:0] mesh_1_7_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177868.4]
  wire [18:0] mesh_1_7_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177868.4]
  wire [(dbits-1):0] mesh_1_7_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177868.4]
  wire  mesh_1_7_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177868.4]
  wire [5:0] mesh_1_7_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177868.4]
  wire [7:0] mesh_1_7_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177868.4]
  wire [(dbits-1):0] mesh_1_7_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177868.4]
  wire [18:0] mesh_1_7_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177868.4]
  wire  mesh_1_7_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177868.4]
  wire [5:0] mesh_1_7_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177868.4]
  wire  mesh_1_7_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177868.4]
  wire  mesh_1_7_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177868.4]
  wire  mesh_2_0_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177871.4]
  wire [7:0] mesh_2_0_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177871.4]
  wire [18:0] mesh_2_0_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177871.4]
  wire [(dbits-1):0] mesh_2_0_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177871.4]
  wire  mesh_2_0_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177871.4]
  wire [5:0] mesh_2_0_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177871.4]
  wire [7:0] mesh_2_0_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177871.4]
  wire [(dbits-1):0] mesh_2_0_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177871.4]
  wire [18:0] mesh_2_0_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177871.4]
  wire  mesh_2_0_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177871.4]
  wire [5:0] mesh_2_0_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177871.4]
  wire  mesh_2_0_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177871.4]
  wire  mesh_2_0_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177871.4]
  wire  mesh_2_1_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177874.4]
  wire [7:0] mesh_2_1_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177874.4]
  wire [18:0] mesh_2_1_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177874.4]
  wire [(dbits-1):0] mesh_2_1_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177874.4]
  wire  mesh_2_1_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177874.4]
  wire [5:0] mesh_2_1_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177874.4]
  wire [7:0] mesh_2_1_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177874.4]
  wire [(dbits-1):0] mesh_2_1_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177874.4]
  wire [18:0] mesh_2_1_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177874.4]
  wire  mesh_2_1_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177874.4]
  wire [5:0] mesh_2_1_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177874.4]
  wire  mesh_2_1_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177874.4]
  wire  mesh_2_1_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177874.4]
  wire  mesh_2_2_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177877.4]
  wire [7:0] mesh_2_2_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177877.4]
  wire [18:0] mesh_2_2_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177877.4]
  wire [(dbits-1):0] mesh_2_2_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177877.4]
  wire  mesh_2_2_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177877.4]
  wire [5:0] mesh_2_2_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177877.4]
  wire [7:0] mesh_2_2_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177877.4]
  wire [(dbits-1):0] mesh_2_2_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177877.4]
  wire [18:0] mesh_2_2_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177877.4]
  wire  mesh_2_2_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177877.4]
  wire [5:0] mesh_2_2_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177877.4]
  wire  mesh_2_2_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177877.4]
  wire  mesh_2_2_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177877.4]
  wire  mesh_2_3_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177880.4]
  wire [7:0] mesh_2_3_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177880.4]
  wire [18:0] mesh_2_3_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177880.4]
  wire [(dbits-1):0] mesh_2_3_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177880.4]
  wire  mesh_2_3_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177880.4]
  wire [5:0] mesh_2_3_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177880.4]
  wire [7:0] mesh_2_3_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177880.4]
  wire [(dbits-1):0] mesh_2_3_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177880.4]
  wire [18:0] mesh_2_3_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177880.4]
  wire  mesh_2_3_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177880.4]
  wire [5:0] mesh_2_3_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177880.4]
  wire  mesh_2_3_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177880.4]
  wire  mesh_2_3_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177880.4]
  wire  mesh_2_4_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177883.4]
  wire [7:0] mesh_2_4_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177883.4]
  wire [18:0] mesh_2_4_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177883.4]
  wire [(dbits-1):0] mesh_2_4_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177883.4]
  wire  mesh_2_4_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177883.4]
  wire [5:0] mesh_2_4_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177883.4]
  wire [7:0] mesh_2_4_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177883.4]
  wire [(dbits-1):0] mesh_2_4_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177883.4]
  wire [18:0] mesh_2_4_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177883.4]
  wire  mesh_2_4_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177883.4]
  wire [5:0] mesh_2_4_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177883.4]
  wire  mesh_2_4_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177883.4]
  wire  mesh_2_4_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177883.4]
  wire  mesh_2_5_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177886.4]
  wire [7:0] mesh_2_5_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177886.4]
  wire [18:0] mesh_2_5_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177886.4]
  wire [(dbits-1):0] mesh_2_5_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177886.4]
  wire  mesh_2_5_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177886.4]
  wire [5:0] mesh_2_5_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177886.4]
  wire [7:0] mesh_2_5_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177886.4]
  wire [(dbits-1):0] mesh_2_5_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177886.4]
  wire [18:0] mesh_2_5_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177886.4]
  wire  mesh_2_5_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177886.4]
  wire [5:0] mesh_2_5_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177886.4]
  wire  mesh_2_5_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177886.4]
  wire  mesh_2_5_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177886.4]
  wire  mesh_2_6_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177889.4]
  wire [7:0] mesh_2_6_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177889.4]
  wire [18:0] mesh_2_6_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177889.4]
  wire [(dbits-1):0] mesh_2_6_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177889.4]
  wire  mesh_2_6_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177889.4]
  wire [5:0] mesh_2_6_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177889.4]
  wire [7:0] mesh_2_6_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177889.4]
  wire [(dbits-1):0] mesh_2_6_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177889.4]
  wire [18:0] mesh_2_6_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177889.4]
  wire  mesh_2_6_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177889.4]
  wire [5:0] mesh_2_6_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177889.4]
  wire  mesh_2_6_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177889.4]
  wire  mesh_2_6_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177889.4]
  wire  mesh_2_7_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177892.4]
  wire [7:0] mesh_2_7_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177892.4]
  wire [18:0] mesh_2_7_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177892.4]
  wire [(dbits-1):0] mesh_2_7_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177892.4]
  wire  mesh_2_7_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177892.4]
  wire [5:0] mesh_2_7_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177892.4]
  wire [7:0] mesh_2_7_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177892.4]
  wire [(dbits-1):0] mesh_2_7_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177892.4]
  wire [18:0] mesh_2_7_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177892.4]
  wire  mesh_2_7_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177892.4]
  wire [5:0] mesh_2_7_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177892.4]
  wire  mesh_2_7_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177892.4]
  wire  mesh_2_7_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177892.4]
  wire  mesh_3_0_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177895.4]
  wire [7:0] mesh_3_0_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177895.4]
  wire [18:0] mesh_3_0_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177895.4]
  wire [(dbits-1):0] mesh_3_0_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177895.4]
  wire  mesh_3_0_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177895.4]
  wire [5:0] mesh_3_0_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177895.4]
  wire [7:0] mesh_3_0_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177895.4]
  wire [(dbits-1):0] mesh_3_0_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177895.4]
  wire [18:0] mesh_3_0_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177895.4]
  wire  mesh_3_0_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177895.4]
  wire [5:0] mesh_3_0_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177895.4]
  wire  mesh_3_0_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177895.4]
  wire  mesh_3_0_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177895.4]
  wire  mesh_3_1_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177898.4]
  wire [7:0] mesh_3_1_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177898.4]
  wire [18:0] mesh_3_1_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177898.4]
  wire [(dbits-1):0] mesh_3_1_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177898.4]
  wire  mesh_3_1_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177898.4]
  wire [5:0] mesh_3_1_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177898.4]
  wire [7:0] mesh_3_1_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177898.4]
  wire [(dbits-1):0] mesh_3_1_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177898.4]
  wire [18:0] mesh_3_1_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177898.4]
  wire  mesh_3_1_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177898.4]
  wire [5:0] mesh_3_1_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177898.4]
  wire  mesh_3_1_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177898.4]
  wire  mesh_3_1_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177898.4]
  wire  mesh_3_2_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177901.4]
  wire [7:0] mesh_3_2_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177901.4]
  wire [18:0] mesh_3_2_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177901.4]
  wire [(dbits-1):0] mesh_3_2_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177901.4]
  wire  mesh_3_2_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177901.4]
  wire [5:0] mesh_3_2_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177901.4]
  wire [7:0] mesh_3_2_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177901.4]
  wire [(dbits-1):0] mesh_3_2_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177901.4]
  wire [18:0] mesh_3_2_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177901.4]
  wire  mesh_3_2_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177901.4]
  wire [5:0] mesh_3_2_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177901.4]
  wire  mesh_3_2_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177901.4]
  wire  mesh_3_2_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177901.4]
  wire  mesh_3_3_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177904.4]
  wire [7:0] mesh_3_3_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177904.4]
  wire [18:0] mesh_3_3_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177904.4]
  wire [(dbits-1):0] mesh_3_3_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177904.4]
  wire  mesh_3_3_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177904.4]
  wire [5:0] mesh_3_3_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177904.4]
  wire [7:0] mesh_3_3_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177904.4]
  wire [(dbits-1):0] mesh_3_3_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177904.4]
  wire [18:0] mesh_3_3_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177904.4]
  wire  mesh_3_3_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177904.4]
  wire [5:0] mesh_3_3_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177904.4]
  wire  mesh_3_3_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177904.4]
  wire  mesh_3_3_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177904.4]
  wire  mesh_3_4_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177907.4]
  wire [7:0] mesh_3_4_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177907.4]
  wire [18:0] mesh_3_4_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177907.4]
  wire [(dbits-1):0] mesh_3_4_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177907.4]
  wire  mesh_3_4_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177907.4]
  wire [5:0] mesh_3_4_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177907.4]
  wire [7:0] mesh_3_4_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177907.4]
  wire [(dbits-1):0] mesh_3_4_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177907.4]
  wire [18:0] mesh_3_4_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177907.4]
  wire  mesh_3_4_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177907.4]
  wire [5:0] mesh_3_4_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177907.4]
  wire  mesh_3_4_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177907.4]
  wire  mesh_3_4_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177907.4]
  wire  mesh_3_5_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177910.4]
  wire [7:0] mesh_3_5_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177910.4]
  wire [18:0] mesh_3_5_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177910.4]
  wire [(dbits-1):0] mesh_3_5_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177910.4]
  wire  mesh_3_5_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177910.4]
  wire [5:0] mesh_3_5_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177910.4]
  wire [7:0] mesh_3_5_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177910.4]
  wire [(dbits-1):0] mesh_3_5_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177910.4]
  wire [18:0] mesh_3_5_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177910.4]
  wire  mesh_3_5_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177910.4]
  wire [5:0] mesh_3_5_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177910.4]
  wire  mesh_3_5_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177910.4]
  wire  mesh_3_5_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177910.4]
  wire  mesh_3_6_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177913.4]
  wire [7:0] mesh_3_6_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177913.4]
  wire [18:0] mesh_3_6_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177913.4]
  wire [(dbits-1):0] mesh_3_6_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177913.4]
  wire  mesh_3_6_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177913.4]
  wire [5:0] mesh_3_6_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177913.4]
  wire [7:0] mesh_3_6_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177913.4]
  wire [(dbits-1):0] mesh_3_6_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177913.4]
  wire [18:0] mesh_3_6_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177913.4]
  wire  mesh_3_6_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177913.4]
  wire [5:0] mesh_3_6_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177913.4]
  wire  mesh_3_6_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177913.4]
  wire  mesh_3_6_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177913.4]
  wire  mesh_3_7_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177916.4]
  wire [7:0] mesh_3_7_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177916.4]
  wire [18:0] mesh_3_7_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177916.4]
  wire [(dbits-1):0] mesh_3_7_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177916.4]
  wire  mesh_3_7_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177916.4]
  wire [5:0] mesh_3_7_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177916.4]
  wire [7:0] mesh_3_7_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177916.4]
  wire [(dbits-1):0] mesh_3_7_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177916.4]
  wire [18:0] mesh_3_7_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177916.4]
  wire  mesh_3_7_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177916.4]
  wire [5:0] mesh_3_7_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177916.4]
  wire  mesh_3_7_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177916.4]
  wire  mesh_3_7_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177916.4]
  wire  mesh_4_0_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177919.4]
  wire [7:0] mesh_4_0_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177919.4]
  wire [18:0] mesh_4_0_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177919.4]
  wire [(dbits-1):0] mesh_4_0_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177919.4]
  wire  mesh_4_0_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177919.4]
  wire [5:0] mesh_4_0_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177919.4]
  wire [7:0] mesh_4_0_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177919.4]
  wire [(dbits-1):0] mesh_4_0_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177919.4]
  wire [18:0] mesh_4_0_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177919.4]
  wire  mesh_4_0_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177919.4]
  wire [5:0] mesh_4_0_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177919.4]
  wire  mesh_4_0_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177919.4]
  wire  mesh_4_0_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177919.4]
  wire  mesh_4_1_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177922.4]
  wire [7:0] mesh_4_1_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177922.4]
  wire [18:0] mesh_4_1_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177922.4]
  wire [(dbits-1):0] mesh_4_1_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177922.4]
  wire  mesh_4_1_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177922.4]
  wire [5:0] mesh_4_1_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177922.4]
  wire [7:0] mesh_4_1_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177922.4]
  wire [(dbits-1):0] mesh_4_1_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177922.4]
  wire [18:0] mesh_4_1_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177922.4]
  wire  mesh_4_1_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177922.4]
  wire [5:0] mesh_4_1_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177922.4]
  wire  mesh_4_1_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177922.4]
  wire  mesh_4_1_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177922.4]
  wire  mesh_4_2_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177925.4]
  wire [7:0] mesh_4_2_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177925.4]
  wire [18:0] mesh_4_2_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177925.4]
  wire [(dbits-1):0] mesh_4_2_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177925.4]
  wire  mesh_4_2_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177925.4]
  wire [5:0] mesh_4_2_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177925.4]
  wire [7:0] mesh_4_2_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177925.4]
  wire [(dbits-1):0] mesh_4_2_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177925.4]
  wire [18:0] mesh_4_2_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177925.4]
  wire  mesh_4_2_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177925.4]
  wire [5:0] mesh_4_2_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177925.4]
  wire  mesh_4_2_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177925.4]
  wire  mesh_4_2_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177925.4]
  wire  mesh_4_3_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177928.4]
  wire [7:0] mesh_4_3_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177928.4]
  wire [18:0] mesh_4_3_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177928.4]
  wire [(dbits-1):0] mesh_4_3_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177928.4]
  wire  mesh_4_3_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177928.4]
  wire [5:0] mesh_4_3_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177928.4]
  wire [7:0] mesh_4_3_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177928.4]
  wire [(dbits-1):0] mesh_4_3_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177928.4]
  wire [18:0] mesh_4_3_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177928.4]
  wire  mesh_4_3_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177928.4]
  wire [5:0] mesh_4_3_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177928.4]
  wire  mesh_4_3_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177928.4]
  wire  mesh_4_3_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177928.4]
  wire  mesh_4_4_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177931.4]
  wire [7:0] mesh_4_4_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177931.4]
  wire [18:0] mesh_4_4_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177931.4]
  wire [(dbits-1):0] mesh_4_4_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177931.4]
  wire  mesh_4_4_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177931.4]
  wire [5:0] mesh_4_4_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177931.4]
  wire [7:0] mesh_4_4_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177931.4]
  wire [(dbits-1):0] mesh_4_4_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177931.4]
  wire [18:0] mesh_4_4_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177931.4]
  wire  mesh_4_4_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177931.4]
  wire [5:0] mesh_4_4_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177931.4]
  wire  mesh_4_4_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177931.4]
  wire  mesh_4_4_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177931.4]
  wire  mesh_4_5_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177934.4]
  wire [7:0] mesh_4_5_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177934.4]
  wire [18:0] mesh_4_5_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177934.4]
  wire [(dbits-1):0] mesh_4_5_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177934.4]
  wire  mesh_4_5_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177934.4]
  wire [5:0] mesh_4_5_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177934.4]
  wire [7:0] mesh_4_5_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177934.4]
  wire [(dbits-1):0] mesh_4_5_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177934.4]
  wire [18:0] mesh_4_5_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177934.4]
  wire  mesh_4_5_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177934.4]
  wire [5:0] mesh_4_5_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177934.4]
  wire  mesh_4_5_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177934.4]
  wire  mesh_4_5_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177934.4]
  wire  mesh_4_6_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177937.4]
  wire [7:0] mesh_4_6_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177937.4]
  wire [18:0] mesh_4_6_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177937.4]
  wire [(dbits-1):0] mesh_4_6_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177937.4]
  wire  mesh_4_6_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177937.4]
  wire [5:0] mesh_4_6_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177937.4]
  wire [7:0] mesh_4_6_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177937.4]
  wire [(dbits-1):0] mesh_4_6_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177937.4]
  wire [18:0] mesh_4_6_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177937.4]
  wire  mesh_4_6_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177937.4]
  wire [5:0] mesh_4_6_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177937.4]
  wire  mesh_4_6_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177937.4]
  wire  mesh_4_6_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177937.4]
  wire  mesh_4_7_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177940.4]
  wire [7:0] mesh_4_7_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177940.4]
  wire [18:0] mesh_4_7_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177940.4]
  wire [(dbits-1):0] mesh_4_7_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177940.4]
  wire  mesh_4_7_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177940.4]
  wire [5:0] mesh_4_7_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177940.4]
  wire [7:0] mesh_4_7_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177940.4]
  wire [(dbits-1):0] mesh_4_7_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177940.4]
  wire [18:0] mesh_4_7_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177940.4]
  wire  mesh_4_7_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177940.4]
  wire [5:0] mesh_4_7_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177940.4]
  wire  mesh_4_7_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177940.4]
  wire  mesh_4_7_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177940.4]
  wire  mesh_5_0_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177943.4]
  wire [7:0] mesh_5_0_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177943.4]
  wire [18:0] mesh_5_0_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177943.4]
  wire [(dbits-1):0] mesh_5_0_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177943.4]
  wire  mesh_5_0_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177943.4]
  wire [5:0] mesh_5_0_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177943.4]
  wire [7:0] mesh_5_0_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177943.4]
  wire [(dbits-1):0] mesh_5_0_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177943.4]
  wire [18:0] mesh_5_0_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177943.4]
  wire  mesh_5_0_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177943.4]
  wire [5:0] mesh_5_0_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177943.4]
  wire  mesh_5_0_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177943.4]
  wire  mesh_5_0_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177943.4]
  wire  mesh_5_1_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177946.4]
  wire [7:0] mesh_5_1_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177946.4]
  wire [18:0] mesh_5_1_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177946.4]
  wire [(dbits-1):0] mesh_5_1_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177946.4]
  wire  mesh_5_1_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177946.4]
  wire [5:0] mesh_5_1_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177946.4]
  wire [7:0] mesh_5_1_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177946.4]
  wire [(dbits-1):0] mesh_5_1_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177946.4]
  wire [18:0] mesh_5_1_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177946.4]
  wire  mesh_5_1_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177946.4]
  wire [5:0] mesh_5_1_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177946.4]
  wire  mesh_5_1_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177946.4]
  wire  mesh_5_1_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177946.4]
  wire  mesh_5_2_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177949.4]
  wire [7:0] mesh_5_2_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177949.4]
  wire [18:0] mesh_5_2_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177949.4]
  wire [(dbits-1):0] mesh_5_2_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177949.4]
  wire  mesh_5_2_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177949.4]
  wire [5:0] mesh_5_2_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177949.4]
  wire [7:0] mesh_5_2_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177949.4]
  wire [(dbits-1):0] mesh_5_2_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177949.4]
  wire [18:0] mesh_5_2_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177949.4]
  wire  mesh_5_2_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177949.4]
  wire [5:0] mesh_5_2_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177949.4]
  wire  mesh_5_2_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177949.4]
  wire  mesh_5_2_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177949.4]
  wire  mesh_5_3_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177952.4]
  wire [7:0] mesh_5_3_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177952.4]
  wire [18:0] mesh_5_3_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177952.4]
  wire [(dbits-1):0] mesh_5_3_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177952.4]
  wire  mesh_5_3_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177952.4]
  wire [5:0] mesh_5_3_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177952.4]
  wire [7:0] mesh_5_3_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177952.4]
  wire [(dbits-1):0] mesh_5_3_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177952.4]
  wire [18:0] mesh_5_3_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177952.4]
  wire  mesh_5_3_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177952.4]
  wire [5:0] mesh_5_3_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177952.4]
  wire  mesh_5_3_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177952.4]
  wire  mesh_5_3_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177952.4]
  wire  mesh_5_4_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177955.4]
  wire [7:0] mesh_5_4_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177955.4]
  wire [18:0] mesh_5_4_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177955.4]
  wire [(dbits-1):0] mesh_5_4_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177955.4]
  wire  mesh_5_4_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177955.4]
  wire [5:0] mesh_5_4_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177955.4]
  wire [7:0] mesh_5_4_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177955.4]
  wire [(dbits-1):0] mesh_5_4_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177955.4]
  wire [18:0] mesh_5_4_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177955.4]
  wire  mesh_5_4_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177955.4]
  wire [5:0] mesh_5_4_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177955.4]
  wire  mesh_5_4_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177955.4]
  wire  mesh_5_4_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177955.4]
  wire  mesh_5_5_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177958.4]
  wire [7:0] mesh_5_5_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177958.4]
  wire [18:0] mesh_5_5_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177958.4]
  wire [(dbits-1):0] mesh_5_5_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177958.4]
  wire  mesh_5_5_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177958.4]
  wire [5:0] mesh_5_5_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177958.4]
  wire [7:0] mesh_5_5_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177958.4]
  wire [(dbits-1):0] mesh_5_5_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177958.4]
  wire [18:0] mesh_5_5_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177958.4]
  wire  mesh_5_5_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177958.4]
  wire [5:0] mesh_5_5_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177958.4]
  wire  mesh_5_5_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177958.4]
  wire  mesh_5_5_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177958.4]
  wire  mesh_5_6_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177961.4]
  wire [7:0] mesh_5_6_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177961.4]
  wire [18:0] mesh_5_6_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177961.4]
  wire [(dbits-1):0] mesh_5_6_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177961.4]
  wire  mesh_5_6_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177961.4]
  wire [5:0] mesh_5_6_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177961.4]
  wire [7:0] mesh_5_6_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177961.4]
  wire [(dbits-1):0] mesh_5_6_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177961.4]
  wire [18:0] mesh_5_6_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177961.4]
  wire  mesh_5_6_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177961.4]
  wire [5:0] mesh_5_6_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177961.4]
  wire  mesh_5_6_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177961.4]
  wire  mesh_5_6_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177961.4]
  wire  mesh_5_7_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177964.4]
  wire [7:0] mesh_5_7_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177964.4]
  wire [18:0] mesh_5_7_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177964.4]
  wire [(dbits-1):0] mesh_5_7_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177964.4]
  wire  mesh_5_7_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177964.4]
  wire [5:0] mesh_5_7_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177964.4]
  wire [7:0] mesh_5_7_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177964.4]
  wire [(dbits-1):0] mesh_5_7_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177964.4]
  wire [18:0] mesh_5_7_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177964.4]
  wire  mesh_5_7_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177964.4]
  wire [5:0] mesh_5_7_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177964.4]
  wire  mesh_5_7_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177964.4]
  wire  mesh_5_7_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177964.4]
  wire  mesh_6_0_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177967.4]
  wire [7:0] mesh_6_0_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177967.4]
  wire [18:0] mesh_6_0_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177967.4]
  wire [(dbits-1):0] mesh_6_0_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177967.4]
  wire  mesh_6_0_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177967.4]
  wire [5:0] mesh_6_0_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177967.4]
  wire [7:0] mesh_6_0_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177967.4]
  wire [(dbits-1):0] mesh_6_0_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177967.4]
  wire [18:0] mesh_6_0_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177967.4]
  wire  mesh_6_0_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177967.4]
  wire [5:0] mesh_6_0_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177967.4]
  wire  mesh_6_0_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177967.4]
  wire  mesh_6_0_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177967.4]
  wire  mesh_6_1_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177970.4]
  wire [7:0] mesh_6_1_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177970.4]
  wire [18:0] mesh_6_1_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177970.4]
  wire [(dbits-1):0] mesh_6_1_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177970.4]
  wire  mesh_6_1_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177970.4]
  wire [5:0] mesh_6_1_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177970.4]
  wire [7:0] mesh_6_1_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177970.4]
  wire [(dbits-1):0] mesh_6_1_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177970.4]
  wire [18:0] mesh_6_1_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177970.4]
  wire  mesh_6_1_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177970.4]
  wire [5:0] mesh_6_1_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177970.4]
  wire  mesh_6_1_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177970.4]
  wire  mesh_6_1_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177970.4]
  wire  mesh_6_2_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177973.4]
  wire [7:0] mesh_6_2_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177973.4]
  wire [18:0] mesh_6_2_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177973.4]
  wire [(dbits-1):0] mesh_6_2_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177973.4]
  wire  mesh_6_2_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177973.4]
  wire [5:0] mesh_6_2_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177973.4]
  wire [7:0] mesh_6_2_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177973.4]
  wire [(dbits-1):0] mesh_6_2_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177973.4]
  wire [18:0] mesh_6_2_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177973.4]
  wire  mesh_6_2_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177973.4]
  wire [5:0] mesh_6_2_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177973.4]
  wire  mesh_6_2_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177973.4]
  wire  mesh_6_2_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177973.4]
  wire  mesh_6_3_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177976.4]
  wire [7:0] mesh_6_3_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177976.4]
  wire [18:0] mesh_6_3_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177976.4]
  wire [(dbits-1):0] mesh_6_3_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177976.4]
  wire  mesh_6_3_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177976.4]
  wire [5:0] mesh_6_3_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177976.4]
  wire [7:0] mesh_6_3_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177976.4]
  wire [(dbits-1):0] mesh_6_3_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177976.4]
  wire [18:0] mesh_6_3_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177976.4]
  wire  mesh_6_3_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177976.4]
  wire [5:0] mesh_6_3_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177976.4]
  wire  mesh_6_3_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177976.4]
  wire  mesh_6_3_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177976.4]
  wire  mesh_6_4_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177979.4]
  wire [7:0] mesh_6_4_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177979.4]
  wire [18:0] mesh_6_4_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177979.4]
  wire [(dbits-1):0] mesh_6_4_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177979.4]
  wire  mesh_6_4_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177979.4]
  wire [5:0] mesh_6_4_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177979.4]
  wire [7:0] mesh_6_4_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177979.4]
  wire [(dbits-1):0] mesh_6_4_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177979.4]
  wire [18:0] mesh_6_4_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177979.4]
  wire  mesh_6_4_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177979.4]
  wire [5:0] mesh_6_4_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177979.4]
  wire  mesh_6_4_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177979.4]
  wire  mesh_6_4_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177979.4]
  wire  mesh_6_5_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177982.4]
  wire [7:0] mesh_6_5_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177982.4]
  wire [18:0] mesh_6_5_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177982.4]
  wire [(dbits-1):0] mesh_6_5_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177982.4]
  wire  mesh_6_5_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177982.4]
  wire [5:0] mesh_6_5_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177982.4]
  wire [7:0] mesh_6_5_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177982.4]
  wire [(dbits-1):0] mesh_6_5_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177982.4]
  wire [18:0] mesh_6_5_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177982.4]
  wire  mesh_6_5_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177982.4]
  wire [5:0] mesh_6_5_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177982.4]
  wire  mesh_6_5_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177982.4]
  wire  mesh_6_5_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177982.4]
  wire  mesh_6_6_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177985.4]
  wire [7:0] mesh_6_6_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177985.4]
  wire [18:0] mesh_6_6_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177985.4]
  wire [(dbits-1):0] mesh_6_6_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177985.4]
  wire  mesh_6_6_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177985.4]
  wire [5:0] mesh_6_6_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177985.4]
  wire [7:0] mesh_6_6_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177985.4]
  wire [(dbits-1):0] mesh_6_6_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177985.4]
  wire [18:0] mesh_6_6_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177985.4]
  wire  mesh_6_6_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177985.4]
  wire [5:0] mesh_6_6_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177985.4]
  wire  mesh_6_6_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177985.4]
  wire  mesh_6_6_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177985.4]
  wire  mesh_6_7_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177988.4]
  wire [7:0] mesh_6_7_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177988.4]
  wire [18:0] mesh_6_7_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177988.4]
  wire [(dbits-1):0] mesh_6_7_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177988.4]
  wire  mesh_6_7_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177988.4]
  wire [5:0] mesh_6_7_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177988.4]
  wire [7:0] mesh_6_7_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177988.4]
  wire [(dbits-1):0] mesh_6_7_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177988.4]
  wire [18:0] mesh_6_7_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177988.4]
  wire  mesh_6_7_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177988.4]
  wire [5:0] mesh_6_7_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177988.4]
  wire  mesh_6_7_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177988.4]
  wire  mesh_6_7_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177988.4]
  wire  mesh_7_0_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177991.4]
  wire [7:0] mesh_7_0_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177991.4]
  wire [18:0] mesh_7_0_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177991.4]
  wire [(dbits-1):0] mesh_7_0_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177991.4]
  wire  mesh_7_0_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177991.4]
  wire [5:0] mesh_7_0_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177991.4]
  wire [7:0] mesh_7_0_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177991.4]
  wire [(dbits-1):0] mesh_7_0_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177991.4]
  wire [18:0] mesh_7_0_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177991.4]
  wire  mesh_7_0_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177991.4]
  wire [5:0] mesh_7_0_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177991.4]
  wire  mesh_7_0_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177991.4]
  wire  mesh_7_0_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177991.4]
  wire  mesh_7_1_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177994.4]
  wire [7:0] mesh_7_1_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177994.4]
  wire [18:0] mesh_7_1_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177994.4]
  wire [(dbits-1):0] mesh_7_1_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177994.4]
  wire  mesh_7_1_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177994.4]
  wire [5:0] mesh_7_1_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177994.4]
  wire [7:0] mesh_7_1_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177994.4]
  wire [(dbits-1):0] mesh_7_1_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177994.4]
  wire [18:0] mesh_7_1_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177994.4]
  wire  mesh_7_1_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177994.4]
  wire [5:0] mesh_7_1_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177994.4]
  wire  mesh_7_1_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177994.4]
  wire  mesh_7_1_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177994.4]
  wire  mesh_7_2_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177997.4]
  wire [7:0] mesh_7_2_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177997.4]
  wire [18:0] mesh_7_2_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177997.4]
  wire [(dbits-1):0] mesh_7_2_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177997.4]
  wire  mesh_7_2_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177997.4]
  wire [5:0] mesh_7_2_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177997.4]
  wire [7:0] mesh_7_2_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177997.4]
  wire [(dbits-1):0] mesh_7_2_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177997.4]
  wire [18:0] mesh_7_2_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177997.4]
  wire  mesh_7_2_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177997.4]
  wire [5:0] mesh_7_2_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177997.4]
  wire  mesh_7_2_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177997.4]
  wire  mesh_7_2_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177997.4]
  wire  mesh_7_3_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178000.4]
  wire [7:0] mesh_7_3_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178000.4]
  wire [18:0] mesh_7_3_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178000.4]
  wire [(dbits-1):0] mesh_7_3_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178000.4]
  wire  mesh_7_3_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178000.4]
  wire [5:0] mesh_7_3_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178000.4]
  wire [7:0] mesh_7_3_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178000.4]
  wire [(dbits-1):0] mesh_7_3_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178000.4]
  wire [18:0] mesh_7_3_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178000.4]
  wire  mesh_7_3_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178000.4]
  wire [5:0] mesh_7_3_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178000.4]
  wire  mesh_7_3_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178000.4]
  wire  mesh_7_3_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178000.4]
  wire  mesh_7_4_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178003.4]
  wire [7:0] mesh_7_4_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178003.4]
  wire [18:0] mesh_7_4_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178003.4]
  wire [(dbits-1):0] mesh_7_4_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178003.4]
  wire  mesh_7_4_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178003.4]
  wire [5:0] mesh_7_4_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178003.4]
  wire [7:0] mesh_7_4_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178003.4]
  wire [(dbits-1):0] mesh_7_4_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178003.4]
  wire [18:0] mesh_7_4_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178003.4]
  wire  mesh_7_4_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178003.4]
  wire [5:0] mesh_7_4_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178003.4]
  wire  mesh_7_4_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178003.4]
  wire  mesh_7_4_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178003.4]
  wire  mesh_7_5_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178006.4]
  wire [7:0] mesh_7_5_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178006.4]
  wire [18:0] mesh_7_5_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178006.4]
  wire [(dbits-1):0] mesh_7_5_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178006.4]
  wire  mesh_7_5_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178006.4]
  wire [5:0] mesh_7_5_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178006.4]
  wire [7:0] mesh_7_5_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178006.4]
  wire [(dbits-1):0] mesh_7_5_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178006.4]
  wire [18:0] mesh_7_5_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178006.4]
  wire  mesh_7_5_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178006.4]
  wire [5:0] mesh_7_5_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178006.4]
  wire  mesh_7_5_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178006.4]
  wire  mesh_7_5_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178006.4]
  wire  mesh_7_6_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178009.4]
  wire [7:0] mesh_7_6_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178009.4]
  wire [18:0] mesh_7_6_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178009.4]
  wire [(dbits-1):0] mesh_7_6_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178009.4]
  wire  mesh_7_6_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178009.4]
  wire [5:0] mesh_7_6_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178009.4]
  wire [7:0] mesh_7_6_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178009.4]
  wire [(dbits-1):0] mesh_7_6_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178009.4]
  wire [18:0] mesh_7_6_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178009.4]
  wire  mesh_7_6_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178009.4]
  wire [5:0] mesh_7_6_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178009.4]
  wire  mesh_7_6_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178009.4]
  wire  mesh_7_6_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178009.4]
  wire  mesh_7_7_clock; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178012.4]
  wire [7:0] mesh_7_7_io_in_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178012.4]
  wire [18:0] mesh_7_7_io_in_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178012.4]
  wire [(dbits-1):0] mesh_7_7_io_in_d_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178012.4]
  wire  mesh_7_7_io_in_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178012.4]
  wire [5:0] mesh_7_7_io_in_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178012.4]
  wire [7:0] mesh_7_7_io_out_a_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178012.4]
  wire [(dbits-1):0] mesh_7_7_io_out_c_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178012.4]
  wire [18:0] mesh_7_7_io_out_b_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178012.4]
  wire  mesh_7_7_io_out_control_0_propagate; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178012.4]
  wire [5:0] mesh_7_7_io_out_control_0_shift; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178012.4]
  wire  mesh_7_7_io_in_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178012.4]
  wire  mesh_7_7_io_out_valid_0; // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178012.4]
  reg [7:0] _T_0; // @[Mesh.scala 40:29:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178015.4]
  reg [31:0] _RAND_0;
  reg [7:0] _T_1_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178017.4]
  reg [31:0] _RAND_1;
  reg [7:0] _T_2_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178020.4]
  reg [31:0] _RAND_2;
  reg [7:0] _T_3_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178023.4]
  reg [31:0] _RAND_3;
  reg [7:0] _T_4_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178026.4]
  reg [31:0] _RAND_4;
  reg [7:0] _T_5_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178029.4]
  reg [31:0] _RAND_5;
  reg [7:0] _T_6_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178032.4]
  reg [31:0] _RAND_6;
  reg [7:0] _T_7_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178035.4]
  reg [31:0] _RAND_7;
  reg [7:0] _T_8_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178038.4]
  reg [31:0] _RAND_8;
  reg [7:0] _T_9_0; // @[Mesh.scala 40:29:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178041.4]
  reg [31:0] _RAND_9;
  reg [7:0] _T_10_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178043.4]
  reg [31:0] _RAND_10;
  reg [7:0] _T_11_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178046.4]
  reg [31:0] _RAND_11;
  reg [7:0] _T_12_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178049.4]
  reg [31:0] _RAND_12;
  reg [7:0] _T_13_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178052.4]
  reg [31:0] _RAND_13;
  reg [7:0] _T_14_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178055.4]
  reg [31:0] _RAND_14;
  reg [7:0] _T_15_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178058.4]
  reg [31:0] _RAND_15;
  reg [7:0] _T_16_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178061.4]
  reg [31:0] _RAND_16;
  reg [7:0] _T_17_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178064.4]
  reg [31:0] _RAND_17;
  reg [7:0] _T_18_0; // @[Mesh.scala 40:29:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178067.4]
  reg [31:0] _RAND_18;
  reg [7:0] _T_19_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178069.4]
  reg [31:0] _RAND_19;
  reg [7:0] _T_20_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178072.4]
  reg [31:0] _RAND_20;
  reg [7:0] _T_21_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178075.4]
  reg [31:0] _RAND_21;
  reg [7:0] _T_22_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178078.4]
  reg [31:0] _RAND_22;
  reg [7:0] _T_23_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178081.4]
  reg [31:0] _RAND_23;
  reg [7:0] _T_24_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178084.4]
  reg [31:0] _RAND_24;
  reg [7:0] _T_25_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178087.4]
  reg [31:0] _RAND_25;
  reg [7:0] _T_26_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178090.4]
  reg [31:0] _RAND_26;
  reg [7:0] _T_27_0; // @[Mesh.scala 40:29:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178093.4]
  reg [31:0] _RAND_27;
  reg [7:0] _T_28_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178095.4]
  reg [31:0] _RAND_28;
  reg [7:0] _T_29_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178098.4]
  reg [31:0] _RAND_29;
  reg [7:0] _T_30_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178101.4]
  reg [31:0] _RAND_30;
  reg [7:0] _T_31_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178104.4]
  reg [31:0] _RAND_31;
  reg [7:0] _T_32_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178107.4]
  reg [31:0] _RAND_32;
  reg [7:0] _T_33_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178110.4]
  reg [31:0] _RAND_33;
  reg [7:0] _T_34_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178113.4]
  reg [31:0] _RAND_34;
  reg [7:0] _T_35_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178116.4]
  reg [31:0] _RAND_35;
  reg [7:0] _T_36_0; // @[Mesh.scala 40:29:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178119.4]
  reg [31:0] _RAND_36;
  reg [7:0] _T_37_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178121.4]
  reg [31:0] _RAND_37;
  reg [7:0] _T_38_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178124.4]
  reg [31:0] _RAND_38;
  reg [7:0] _T_39_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178127.4]
  reg [31:0] _RAND_39;
  reg [7:0] _T_40_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178130.4]
  reg [31:0] _RAND_40;
  reg [7:0] _T_41_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178133.4]
  reg [31:0] _RAND_41;
  reg [7:0] _T_42_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178136.4]
  reg [31:0] _RAND_42;
  reg [7:0] _T_43_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178139.4]
  reg [31:0] _RAND_43;
  reg [7:0] _T_44_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178142.4]
  reg [31:0] _RAND_44;
  reg [7:0] _T_45_0; // @[Mesh.scala 40:29:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178145.4]
  reg [31:0] _RAND_45;
  reg [7:0] _T_46_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178147.4]
  reg [31:0] _RAND_46;
  reg [7:0] _T_47_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178150.4]
  reg [31:0] _RAND_47;
  reg [7:0] _T_48_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178153.4]
  reg [31:0] _RAND_48;
  reg [7:0] _T_49_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178156.4]
  reg [31:0] _RAND_49;
  reg [7:0] _T_50_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178159.4]
  reg [31:0] _RAND_50;
  reg [7:0] _T_51_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178162.4]
  reg [31:0] _RAND_51;
  reg [7:0] _T_52_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178165.4]
  reg [31:0] _RAND_52;
  reg [7:0] _T_53_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178168.4]
  reg [31:0] _RAND_53;
  reg [7:0] _T_54_0; // @[Mesh.scala 40:29:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178171.4]
  reg [31:0] _RAND_54;
  reg [7:0] _T_55_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178173.4]
  reg [31:0] _RAND_55;
  reg [7:0] _T_56_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178176.4]
  reg [31:0] _RAND_56;
  reg [7:0] _T_57_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178179.4]
  reg [31:0] _RAND_57;
  reg [7:0] _T_58_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178182.4]
  reg [31:0] _RAND_58;
  reg [7:0] _T_59_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178185.4]
  reg [31:0] _RAND_59;
  reg [7:0] _T_60_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178188.4]
  reg [31:0] _RAND_60;
  reg [7:0] _T_61_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178191.4]
  reg [31:0] _RAND_61;
  reg [7:0] _T_62_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178194.4]
  reg [31:0] _RAND_62;
  reg [7:0] _T_63_0; // @[Mesh.scala 40:29:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178197.4]
  reg [31:0] _RAND_63;
  reg [7:0] _T_64_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178199.4]
  reg [31:0] _RAND_64;
  reg [7:0] _T_65_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178202.4]
  reg [31:0] _RAND_65;
  reg [7:0] _T_66_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178205.4]
  reg [31:0] _RAND_66;
  reg [7:0] _T_67_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178208.4]
  reg [31:0] _RAND_67;
  reg [7:0] _T_68_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178211.4]
  reg [31:0] _RAND_68;
  reg [7:0] _T_69_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178214.4]
  reg [31:0] _RAND_69;
  reg [7:0] _T_70_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178217.4]
  reg [31:0] _RAND_70;
  reg [7:0] _T_71_0; // @[Mesh.scala 42:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178220.4]
  reg [31:0] _RAND_71;
  reg [7:0] _T_72_0; // @[Mesh.scala 48:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178223.4]
  reg [31:0] _RAND_72;
  reg  _T_73_0; // @[Mesh.scala 48:52:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178225.4]
  reg [31:0] _RAND_73;
  reg [7:0] _T_74_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178227.4]
  reg [31:0] _RAND_74;
  reg [18:0] _T_75_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178232.4]
  reg [31:0] _RAND_75;
  reg [18:0] _T_76_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178237.4]
  reg [31:0] _RAND_76;
  reg [18:0] _T_77_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178242.4]
  reg [31:0] _RAND_77;
  reg [18:0] _T_78_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178247.4]
  reg [31:0] _RAND_78;
  reg [18:0] _T_79_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178252.4]
  reg [31:0] _RAND_79;
  reg [18:0] _T_80_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178257.4]
  reg [31:0] _RAND_80;
  reg [18:0] _T_81_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178262.4]
  reg [31:0] _RAND_81;
  reg [7:0] _T_82_0; // @[Mesh.scala 48:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178267.4]
  reg [31:0] _RAND_82;
  reg  _T_83_0; // @[Mesh.scala 48:52:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178269.4]
  reg [31:0] _RAND_83;
  reg [7:0] _T_84_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178271.4]
  reg [31:0] _RAND_84;
  reg [18:0] _T_85_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178276.4]
  reg [31:0] _RAND_85;
  reg [18:0] _T_86_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178281.4]
  reg [31:0] _RAND_86;
  reg [18:0] _T_87_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178286.4]
  reg [31:0] _RAND_87;
  reg [18:0] _T_88_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178291.4]
  reg [31:0] _RAND_88;
  reg [18:0] _T_89_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178296.4]
  reg [31:0] _RAND_89;
  reg [18:0] _T_90_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178301.4]
  reg [31:0] _RAND_90;
  reg [18:0] _T_91_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178306.4]
  reg [31:0] _RAND_91;
  reg [7:0] _T_92_0; // @[Mesh.scala 48:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178311.4]
  reg [31:0] _RAND_92;
  reg  _T_93_0; // @[Mesh.scala 48:52:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178313.4]
  reg [31:0] _RAND_93;
  reg [7:0] _T_94_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178315.4]
  reg [31:0] _RAND_94;
  reg [18:0] _T_95_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178320.4]
  reg [31:0] _RAND_95;
  reg [18:0] _T_96_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178325.4]
  reg [31:0] _RAND_96;
  reg [18:0] _T_97_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178330.4]
  reg [31:0] _RAND_97;
  reg [18:0] _T_98_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178335.4]
  reg [31:0] _RAND_98;
  reg [18:0] _T_99_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178340.4]
  reg [31:0] _RAND_99;
  reg [18:0] _T_100_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178345.4]
  reg [31:0] _RAND_100;
  reg [18:0] _T_101_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178350.4]
  reg [31:0] _RAND_101;
  reg [7:0] _T_102_0; // @[Mesh.scala 48:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178355.4]
  reg [31:0] _RAND_102;
  reg  _T_103_0; // @[Mesh.scala 48:52:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178357.4]
  reg [31:0] _RAND_103;
  reg [7:0] _T_104_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178359.4]
  reg [31:0] _RAND_104;
  reg [18:0] _T_105_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178364.4]
  reg [31:0] _RAND_105;
  reg [18:0] _T_106_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178369.4]
  reg [31:0] _RAND_106;
  reg [18:0] _T_107_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178374.4]
  reg [31:0] _RAND_107;
  reg [18:0] _T_108_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178379.4]
  reg [31:0] _RAND_108;
  reg [18:0] _T_109_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178384.4]
  reg [31:0] _RAND_109;
  reg [18:0] _T_110_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178389.4]
  reg [31:0] _RAND_110;
  reg [18:0] _T_111_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178394.4]
  reg [31:0] _RAND_111;
  reg [7:0] _T_112_0; // @[Mesh.scala 48:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178399.4]
  reg [31:0] _RAND_112;
  reg  _T_113_0; // @[Mesh.scala 48:52:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178401.4]
  reg [31:0] _RAND_113;
  reg [7:0] _T_114_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178403.4]
  reg [31:0] _RAND_114;
  reg [18:0] _T_115_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178408.4]
  reg [31:0] _RAND_115;
  reg [18:0] _T_116_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178413.4]
  reg [31:0] _RAND_116;
  reg [18:0] _T_117_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178418.4]
  reg [31:0] _RAND_117;
  reg [18:0] _T_118_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178423.4]
  reg [31:0] _RAND_118;
  reg [18:0] _T_119_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178428.4]
  reg [31:0] _RAND_119;
  reg [18:0] _T_120_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178433.4]
  reg [31:0] _RAND_120;
  reg [18:0] _T_121_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178438.4]
  reg [31:0] _RAND_121;
  reg [7:0] _T_122_0; // @[Mesh.scala 48:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178443.4]
  reg [31:0] _RAND_122;
  reg  _T_123_0; // @[Mesh.scala 48:52:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178445.4]
  reg [31:0] _RAND_123;
  reg [7:0] _T_124_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178447.4]
  reg [31:0] _RAND_124;
  reg [18:0] _T_125_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178452.4]
  reg [31:0] _RAND_125;
  reg [18:0] _T_126_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178457.4]
  reg [31:0] _RAND_126;
  reg [18:0] _T_127_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178462.4]
  reg [31:0] _RAND_127;
  reg [18:0] _T_128_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178467.4]
  reg [31:0] _RAND_128;
  reg [18:0] _T_129_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178472.4]
  reg [31:0] _RAND_129;
  reg [18:0] _T_130_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178477.4]
  reg [31:0] _RAND_130;
  reg [18:0] _T_131_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178482.4]
  reg [31:0] _RAND_131;
  reg [7:0] _T_132_0; // @[Mesh.scala 48:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178487.4]
  reg [31:0] _RAND_132;
  reg  _T_133_0; // @[Mesh.scala 48:52:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178489.4]
  reg [31:0] _RAND_133;
  reg [7:0] _T_134_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178491.4]
  reg [31:0] _RAND_134;
  reg [18:0] _T_135_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178496.4]
  reg [31:0] _RAND_135;
  reg [18:0] _T_136_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178501.4]
  reg [31:0] _RAND_136;
  reg [18:0] _T_137_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178506.4]
  reg [31:0] _RAND_137;
  reg [18:0] _T_138_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178511.4]
  reg [31:0] _RAND_138;
  reg [18:0] _T_139_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178516.4]
  reg [31:0] _RAND_139;
  reg [18:0] _T_140_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178521.4]
  reg [31:0] _RAND_140;
  reg [18:0] _T_141_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178526.4]
  reg [31:0] _RAND_141;
  reg [7:0] _T_142_0; // @[Mesh.scala 48:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178531.4]
  reg [31:0] _RAND_142;
  reg  _T_143_0; // @[Mesh.scala 48:52:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178533.4]
  reg [31:0] _RAND_143;
  reg [7:0] _T_144_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178535.4]
  reg [31:0] _RAND_144;
  reg [18:0] _T_145_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178540.4]
  reg [31:0] _RAND_145;
  reg [18:0] _T_146_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178545.4]
  reg [31:0] _RAND_146;
  reg [18:0] _T_147_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178550.4]
  reg [31:0] _RAND_147;
  reg [18:0] _T_148_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178555.4]
  reg [31:0] _RAND_148;
  reg [18:0] _T_149_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178560.4]
  reg [31:0] _RAND_149;
  reg [18:0] _T_150_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178565.4]
  reg [31:0] _RAND_150;
  reg [18:0] _T_151_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178570.4]
  reg [31:0] _RAND_151;
  reg [7:0] _T_152_0; // @[Mesh.scala 56:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178575.4]
  reg [31:0] _RAND_152;
  reg  _T_153_0; // @[Mesh.scala 56:52:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178577.4]
  reg [31:0] _RAND_153;
  reg [7:0] _T_154_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178579.4]
  reg [31:0] _RAND_154;
  reg [(dbits-1):0] _T_155_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178584.4]
  reg [(dbits-1):0] _RAND_155;
  reg [(dbits-1):0] _T_156_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178589.4]
  reg [(dbits-1):0] _RAND_156;
  reg [(dbits-1):0] _T_157_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178594.4]
  reg [(dbits-1):0] _RAND_157;
  reg [(dbits-1):0] _T_158_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178599.4]
  reg [(dbits-1):0] _RAND_158;
  reg [(dbits-1):0] _T_159_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178604.4]
  reg [(dbits-1):0] _RAND_159;
  reg [(dbits-1):0] _T_160_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178609.4]
  reg [(dbits-1):0] _RAND_160;
  reg [(dbits-1):0] _T_161_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178614.4]
  reg [(dbits-1):0] _RAND_161;
  reg [7:0] _T_162_0; // @[Mesh.scala 56:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178619.4]
  reg [31:0] _RAND_162;
  reg  _T_163_0; // @[Mesh.scala 56:52:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178621.4]
  reg [31:0] _RAND_163;
  reg [7:0] _T_164_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178623.4]
  reg [31:0] _RAND_164;
  reg [(dbits-1):0] _T_165_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178628.4]
  reg [(dbits-1):0] _RAND_165;
  reg [(dbits-1):0] _T_166_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178633.4]
  reg [(dbits-1):0] _RAND_166;
  reg [(dbits-1):0] _T_167_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178638.4]
  reg [(dbits-1):0] _RAND_167;
  reg [(dbits-1):0] _T_168_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178643.4]
  reg [(dbits-1):0] _RAND_168;
  reg [(dbits-1):0] _T_169_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178648.4]
  reg [(dbits-1):0] _RAND_169;
  reg [(dbits-1):0] _T_170_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178653.4]
  reg [(dbits-1):0] _RAND_170;
  reg [(dbits-1):0] _T_171_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178658.4]
  reg [(dbits-1):0] _RAND_171;
  reg [7:0] _T_172_0; // @[Mesh.scala 56:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178663.4]
  reg [31:0] _RAND_172;
  reg  _T_173_0; // @[Mesh.scala 56:52:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178665.4]
  reg [31:0] _RAND_173;
  reg [7:0] _T_174_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178667.4]
  reg [31:0] _RAND_174;
  reg [(dbits-1):0] _T_175_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178672.4]
  reg [(dbits-1):0] _RAND_175;
  reg [(dbits-1):0] _T_176_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178677.4]
  reg [(dbits-1):0] _RAND_176;
  reg [(dbits-1):0] _T_177_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178682.4]
  reg [(dbits-1):0] _RAND_177;
  reg [(dbits-1):0] _T_178_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178687.4]
  reg [(dbits-1):0] _RAND_178;
  reg [(dbits-1):0] _T_179_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178692.4]
  reg [(dbits-1):0] _RAND_179;
  reg [(dbits-1):0] _T_180_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178697.4]
  reg [(dbits-1):0] _RAND_180;
  reg [(dbits-1):0] _T_181_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178702.4]
  reg [(dbits-1):0] _RAND_181;
  reg [7:0] _T_182_0; // @[Mesh.scala 56:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178707.4]
  reg [31:0] _RAND_182;
  reg  _T_183_0; // @[Mesh.scala 56:52:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178709.4]
  reg [31:0] _RAND_183;
  reg [7:0] _T_184_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178711.4]
  reg [31:0] _RAND_184;
  reg [(dbits-1):0] _T_185_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178716.4]
  reg [(dbits-1):0] _RAND_185;
  reg [(dbits-1):0] _T_186_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178721.4]
  reg [(dbits-1):0] _RAND_186;
  reg [(dbits-1):0] _T_187_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178726.4]
  reg [(dbits-1):0] _RAND_187;
  reg [(dbits-1):0] _T_188_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178731.4]
  reg [(dbits-1):0] _RAND_188;
  reg [(dbits-1):0] _T_189_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178736.4]
  reg [(dbits-1):0] _RAND_189;
  reg [(dbits-1):0] _T_190_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178741.4]
  reg [(dbits-1):0] _RAND_190;
  reg [(dbits-1):0] _T_191_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178746.4]
  reg [(dbits-1):0] _RAND_191;
  reg [7:0] _T_192_0; // @[Mesh.scala 56:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178751.4]
  reg [31:0] _RAND_192;
  reg  _T_193_0; // @[Mesh.scala 56:52:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178753.4]
  reg [31:0] _RAND_193;
  reg [7:0] _T_194_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178755.4]
  reg [31:0] _RAND_194;
  reg [(dbits-1):0] _T_195_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178760.4]
  reg [(dbits-1):0] _RAND_195;
  reg [(dbits-1):0] _T_196_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178765.4]
  reg [(dbits-1):0] _RAND_196;
  reg [(dbits-1):0] _T_197_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178770.4]
  reg [(dbits-1):0] _RAND_197;
  reg [(dbits-1):0] _T_198_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178775.4]
  reg [(dbits-1):0] _RAND_198;
  reg [(dbits-1):0] _T_199_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178780.4]
  reg [(dbits-1):0] _RAND_199;
  reg [(dbits-1):0] _T_200_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178785.4]
  reg [(dbits-1):0] _RAND_200;
  reg [(dbits-1):0] _T_201_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178790.4]
  reg [(dbits-1):0] _RAND_201;
  reg [7:0] _T_202_0; // @[Mesh.scala 56:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178795.4]
  reg [31:0] _RAND_202;
  reg  _T_203_0; // @[Mesh.scala 56:52:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178797.4]
  reg [31:0] _RAND_203;
  reg [7:0] _T_204_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178799.4]
  reg [31:0] _RAND_204;
  reg [(dbits-1):0] _T_205_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178804.4]
  reg [(dbits-1):0] _RAND_205;
  reg [(dbits-1):0] _T_206_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178809.4]
  reg [(dbits-1):0] _RAND_206;
  reg [(dbits-1):0] _T_207_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178814.4]
  reg [(dbits-1):0] _RAND_207;
  reg [(dbits-1):0] _T_208_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178819.4]
  reg [(dbits-1):0] _RAND_208;
  reg [(dbits-1):0] _T_209_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178824.4]
  reg [(dbits-1):0] _RAND_209;
  reg [(dbits-1):0] _T_210_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178829.4]
  reg [(dbits-1):0] _RAND_210;
  reg [(dbits-1):0] _T_211_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178834.4]
  reg [(dbits-1):0] _RAND_211;
  reg [7:0] _T_212_0; // @[Mesh.scala 56:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178839.4]
  reg [31:0] _RAND_212;
  reg  _T_213_0; // @[Mesh.scala 56:52:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178841.4]
  reg [31:0] _RAND_213;
  reg [7:0] _T_214_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178843.4]
  reg [31:0] _RAND_214;
  reg [(dbits-1):0] _T_215_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178848.4]
  reg [(dbits-1):0] _RAND_215;
  reg [(dbits-1):0] _T_216_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178853.4]
  reg [(dbits-1):0] _RAND_216;
  reg [(dbits-1):0] _T_217_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178858.4]
  reg [(dbits-1):0] _RAND_217;
  reg [(dbits-1):0] _T_218_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178863.4]
  reg [(dbits-1):0] _RAND_218;
  reg [(dbits-1):0] _T_219_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178868.4]
  reg [(dbits-1):0] _RAND_219;
  reg [(dbits-1):0] _T_220_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178873.4]
  reg [(dbits-1):0] _RAND_220;
  reg [(dbits-1):0] _T_221_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178878.4]
  reg [(dbits-1):0] _RAND_221;
  reg [7:0] _T_222_0; // @[Mesh.scala 56:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178883.4]
  reg [31:0] _RAND_222;
  reg  _T_223_0; // @[Mesh.scala 56:52:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178885.4]
  reg [31:0] _RAND_223;
  reg [7:0] _T_224_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178887.4]
  reg [31:0] _RAND_224;
  reg [(dbits-1):0] _T_225_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178892.4]
  reg [(dbits-1):0] _RAND_225;
  reg [(dbits-1):0] _T_226_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178897.4]
  reg [(dbits-1):0] _RAND_226;
  reg [(dbits-1):0] _T_227_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178902.4]
  reg [(dbits-1):0] _RAND_227;
  reg [(dbits-1):0] _T_228_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178907.4]
  reg [(dbits-1):0] _RAND_228;
  reg [(dbits-1):0] _T_229_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178912.4]
  reg [(dbits-1):0] _RAND_229;
  reg [(dbits-1):0] _T_230_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178917.4]
  reg [(dbits-1):0] _RAND_230;
  reg [(dbits-1):0] _T_231_0; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178922.4]
  reg [(dbits-1):0] _RAND_231;
  reg  _T_232_0_propagate; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178927.4]
  reg [31:0] _RAND_232;
  reg [5:0] _T_232_0_shift; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178927.4]
  reg [31:0] _RAND_233;
  reg  _T_233_0; // @[Mesh.scala 64:58:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178931.4]
  reg [31:0] _RAND_234;
  reg [5:0] _T_234; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178933.4]
  reg [31:0] _RAND_235;
  reg  _T_236; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178943.4]
  reg [31:0] _RAND_236;
  reg [5:0] _T_237; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178948.4]
  reg [31:0] _RAND_237;
  reg  _T_239; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178958.4]
  reg [31:0] _RAND_238;
  reg [5:0] _T_240; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178963.4]
  reg [31:0] _RAND_239;
  reg  _T_242; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178973.4]
  reg [31:0] _RAND_240;
  reg [5:0] _T_243; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178978.4]
  reg [31:0] _RAND_241;
  reg  _T_245; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178988.4]
  reg [31:0] _RAND_242;
  reg [5:0] _T_246; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178993.4]
  reg [31:0] _RAND_243;
  reg  _T_248; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179003.4]
  reg [31:0] _RAND_244;
  reg [5:0] _T_249; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179008.4]
  reg [31:0] _RAND_245;
  reg  _T_251; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179018.4]
  reg [31:0] _RAND_246;
  reg [5:0] _T_252; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179023.4]
  reg [31:0] _RAND_247;
  reg  _T_254; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179033.4]
  reg [31:0] _RAND_248;
  reg [5:0] _T_255; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179038.4]
  reg [31:0] _RAND_249;
  reg  _T_257; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179048.4]
  reg [31:0] _RAND_250;
  reg  _T_258_0_propagate; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179053.4]
  reg [31:0] _RAND_251;
  reg [5:0] _T_258_0_shift; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179053.4]
  reg [31:0] _RAND_252;
  reg  _T_259_0; // @[Mesh.scala 64:58:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179057.4]
  reg [31:0] _RAND_253;
  reg [5:0] _T_260; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179059.4]
  reg [31:0] _RAND_254;
  reg  _T_262; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179069.4]
  reg [31:0] _RAND_255;
  reg [5:0] _T_263; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179074.4]
  reg [31:0] _RAND_256;
  reg  _T_265; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179084.4]
  reg [31:0] _RAND_257;
  reg [5:0] _T_266; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179089.4]
  reg [31:0] _RAND_258;
  reg  _T_268; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179099.4]
  reg [31:0] _RAND_259;
  reg [5:0] _T_269; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179104.4]
  reg [31:0] _RAND_260;
  reg  _T_271; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179114.4]
  reg [31:0] _RAND_261;
  reg [5:0] _T_272; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179119.4]
  reg [31:0] _RAND_262;
  reg  _T_274; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179129.4]
  reg [31:0] _RAND_263;
  reg [5:0] _T_275; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179134.4]
  reg [31:0] _RAND_264;
  reg  _T_277; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179144.4]
  reg [31:0] _RAND_265;
  reg [5:0] _T_278; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179149.4]
  reg [31:0] _RAND_266;
  reg  _T_280; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179159.4]
  reg [31:0] _RAND_267;
  reg [5:0] _T_281; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179164.4]
  reg [31:0] _RAND_268;
  reg  _T_283; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179174.4]
  reg [31:0] _RAND_269;
  reg  _T_284_0_propagate; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179179.4]
  reg [31:0] _RAND_270;
  reg [5:0] _T_284_0_shift; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179179.4]
  reg [31:0] _RAND_271;
  reg  _T_285_0; // @[Mesh.scala 64:58:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179183.4]
  reg [31:0] _RAND_272;
  reg [5:0] _T_286; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179185.4]
  reg [31:0] _RAND_273;
  reg  _T_288; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179195.4]
  reg [31:0] _RAND_274;
  reg [5:0] _T_289; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179200.4]
  reg [31:0] _RAND_275;
  reg  _T_291; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179210.4]
  reg [31:0] _RAND_276;
  reg [5:0] _T_292; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179215.4]
  reg [31:0] _RAND_277;
  reg  _T_294; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179225.4]
  reg [31:0] _RAND_278;
  reg [5:0] _T_295; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179230.4]
  reg [31:0] _RAND_279;
  reg  _T_297; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179240.4]
  reg [31:0] _RAND_280;
  reg [5:0] _T_298; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179245.4]
  reg [31:0] _RAND_281;
  reg  _T_300; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179255.4]
  reg [31:0] _RAND_282;
  reg [5:0] _T_301; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179260.4]
  reg [31:0] _RAND_283;
  reg  _T_303; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179270.4]
  reg [31:0] _RAND_284;
  reg [5:0] _T_304; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179275.4]
  reg [31:0] _RAND_285;
  reg  _T_306; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179285.4]
  reg [31:0] _RAND_286;
  reg [5:0] _T_307; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179290.4]
  reg [31:0] _RAND_287;
  reg  _T_309; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179300.4]
  reg [31:0] _RAND_288;
  reg  _T_310_0_propagate; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179305.4]
  reg [31:0] _RAND_289;
  reg [5:0] _T_310_0_shift; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179305.4]
  reg [31:0] _RAND_290;
  reg  _T_311_0; // @[Mesh.scala 64:58:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179309.4]
  reg [31:0] _RAND_291;
  reg [5:0] _T_312; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179311.4]
  reg [31:0] _RAND_292;
  reg  _T_314; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179321.4]
  reg [31:0] _RAND_293;
  reg [5:0] _T_315; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179326.4]
  reg [31:0] _RAND_294;
  reg  _T_317; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179336.4]
  reg [31:0] _RAND_295;
  reg [5:0] _T_318; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179341.4]
  reg [31:0] _RAND_296;
  reg  _T_320; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179351.4]
  reg [31:0] _RAND_297;
  reg [5:0] _T_321; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179356.4]
  reg [31:0] _RAND_298;
  reg  _T_323; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179366.4]
  reg [31:0] _RAND_299;
  reg [5:0] _T_324; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179371.4]
  reg [31:0] _RAND_300;
  reg  _T_326; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179381.4]
  reg [31:0] _RAND_301;
  reg [5:0] _T_327; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179386.4]
  reg [31:0] _RAND_302;
  reg  _T_329; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179396.4]
  reg [31:0] _RAND_303;
  reg [5:0] _T_330; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179401.4]
  reg [31:0] _RAND_304;
  reg  _T_332; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179411.4]
  reg [31:0] _RAND_305;
  reg [5:0] _T_333; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179416.4]
  reg [31:0] _RAND_306;
  reg  _T_335; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179426.4]
  reg [31:0] _RAND_307;
  reg  _T_336_0_propagate; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179431.4]
  reg [31:0] _RAND_308;
  reg [5:0] _T_336_0_shift; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179431.4]
  reg [31:0] _RAND_309;
  reg  _T_337_0; // @[Mesh.scala 64:58:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179435.4]
  reg [31:0] _RAND_310;
  reg [5:0] _T_338; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179437.4]
  reg [31:0] _RAND_311;
  reg  _T_340; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179447.4]
  reg [31:0] _RAND_312;
  reg [5:0] _T_341; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179452.4]
  reg [31:0] _RAND_313;
  reg  _T_343; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179462.4]
  reg [31:0] _RAND_314;
  reg [5:0] _T_344; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179467.4]
  reg [31:0] _RAND_315;
  reg  _T_346; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179477.4]
  reg [31:0] _RAND_316;
  reg [5:0] _T_347; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179482.4]
  reg [31:0] _RAND_317;
  reg  _T_349; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179492.4]
  reg [31:0] _RAND_318;
  reg [5:0] _T_350; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179497.4]
  reg [31:0] _RAND_319;
  reg  _T_352; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179507.4]
  reg [31:0] _RAND_320;
  reg [5:0] _T_353; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179512.4]
  reg [31:0] _RAND_321;
  reg  _T_355; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179522.4]
  reg [31:0] _RAND_322;
  reg [5:0] _T_356; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179527.4]
  reg [31:0] _RAND_323;
  reg  _T_358; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179537.4]
  reg [31:0] _RAND_324;
  reg [5:0] _T_359; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179542.4]
  reg [31:0] _RAND_325;
  reg  _T_361; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179552.4]
  reg [31:0] _RAND_326;
  reg  _T_362_0_propagate; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179557.4]
  reg [31:0] _RAND_327;
  reg [5:0] _T_362_0_shift; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179557.4]
  reg [31:0] _RAND_328;
  reg  _T_363_0; // @[Mesh.scala 64:58:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179561.4]
  reg [31:0] _RAND_329;
  reg [5:0] _T_364; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179563.4]
  reg [31:0] _RAND_330;
  reg  _T_366; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179573.4]
  reg [31:0] _RAND_331;
  reg [5:0] _T_367; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179578.4]
  reg [31:0] _RAND_332;
  reg  _T_369; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179588.4]
  reg [31:0] _RAND_333;
  reg [5:0] _T_370; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179593.4]
  reg [31:0] _RAND_334;
  reg  _T_372; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179603.4]
  reg [31:0] _RAND_335;
  reg [5:0] _T_373; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179608.4]
  reg [31:0] _RAND_336;
  reg  _T_375; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179618.4]
  reg [31:0] _RAND_337;
  reg [5:0] _T_376; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179623.4]
  reg [31:0] _RAND_338;
  reg  _T_378; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179633.4]
  reg [31:0] _RAND_339;
  reg [5:0] _T_379; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179638.4]
  reg [31:0] _RAND_340;
  reg  _T_381; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179648.4]
  reg [31:0] _RAND_341;
  reg [5:0] _T_382; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179653.4]
  reg [31:0] _RAND_342;
  reg  _T_384; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179663.4]
  reg [31:0] _RAND_343;
  reg [5:0] _T_385; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179668.4]
  reg [31:0] _RAND_344;
  reg  _T_387; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179678.4]
  reg [31:0] _RAND_345;
  reg  _T_388_0_propagate; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179683.4]
  reg [31:0] _RAND_346;
  reg [5:0] _T_388_0_shift; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179683.4]
  reg [31:0] _RAND_347;
  reg  _T_389_0; // @[Mesh.scala 64:58:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179687.4]
  reg [31:0] _RAND_348;
  reg [5:0] _T_390; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179689.4]
  reg [31:0] _RAND_349;
  reg  _T_392; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179699.4]
  reg [31:0] _RAND_350;
  reg [5:0] _T_393; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179704.4]
  reg [31:0] _RAND_351;
  reg  _T_395; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179714.4]
  reg [31:0] _RAND_352;
  reg [5:0] _T_396; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179719.4]
  reg [31:0] _RAND_353;
  reg  _T_398; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179729.4]
  reg [31:0] _RAND_354;
  reg [5:0] _T_399; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179734.4]
  reg [31:0] _RAND_355;
  reg  _T_401; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179744.4]
  reg [31:0] _RAND_356;
  reg [5:0] _T_402; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179749.4]
  reg [31:0] _RAND_357;
  reg  _T_404; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179759.4]
  reg [31:0] _RAND_358;
  reg [5:0] _T_405; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179764.4]
  reg [31:0] _RAND_359;
  reg  _T_407; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179774.4]
  reg [31:0] _RAND_360;
  reg [5:0] _T_408; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179779.4]
  reg [31:0] _RAND_361;
  reg  _T_410; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179789.4]
  reg [31:0] _RAND_362;
  reg [5:0] _T_411; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179794.4]
  reg [31:0] _RAND_363;
  reg  _T_413; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179804.4]
  reg [31:0] _RAND_364;
  reg  _T_414_0_propagate; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179809.4]
  reg [31:0] _RAND_365;
  reg [5:0] _T_414_0_shift; // @[Mesh.scala 64:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179809.4]
  reg [31:0] _RAND_366;
  reg  _T_415_0; // @[Mesh.scala 64:58:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179813.4]
  reg [31:0] _RAND_367;
  reg [5:0] _T_416; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179815.4]
  reg [31:0] _RAND_368;
  reg  _T_418; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179825.4]
  reg [31:0] _RAND_369;
  reg [5:0] _T_419; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179830.4]
  reg [31:0] _RAND_370;
  reg  _T_421; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179840.4]
  reg [31:0] _RAND_371;
  reg [5:0] _T_422; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179845.4]
  reg [31:0] _RAND_372;
  reg  _T_424; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179855.4]
  reg [31:0] _RAND_373;
  reg [5:0] _T_425; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179860.4]
  reg [31:0] _RAND_374;
  reg  _T_427; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179870.4]
  reg [31:0] _RAND_375;
  reg [5:0] _T_428; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179875.4]
  reg [31:0] _RAND_376;
  reg  _T_430; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179885.4]
  reg [31:0] _RAND_377;
  reg [5:0] _T_431; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179890.4]
  reg [31:0] _RAND_378;
  reg  _T_433; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179900.4]
  reg [31:0] _RAND_379;
  reg [5:0] _T_434; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179905.4]
  reg [31:0] _RAND_380;
  reg  _T_436; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179915.4]
  reg [31:0] _RAND_381;
  reg [5:0] _T_437; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179920.4]
  reg [31:0] _RAND_382;
  reg  _T_439; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179930.4]
  reg [31:0] _RAND_383;
  reg  _T_440_0; // @[Mesh.scala 76:30:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179935.4]
  reg [31:0] _RAND_384;
  reg  _T_441_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179937.4]
  reg [31:0] _RAND_385;
  reg  _T_442_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179940.4]
  reg [31:0] _RAND_386;
  reg  _T_443_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179943.4]
  reg [31:0] _RAND_387;
  reg  _T_444_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179946.4]
  reg [31:0] _RAND_388;
  reg  _T_445_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179949.4]
  reg [31:0] _RAND_389;
  reg  _T_446_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179952.4]
  reg [31:0] _RAND_390;
  reg  _T_447_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179955.4]
  reg [31:0] _RAND_391;
  reg  _T_448_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179958.4]
  reg [31:0] _RAND_392;
  reg  _T_449_0; // @[Mesh.scala 76:30:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179961.4]
  reg [31:0] _RAND_393;
  reg  _T_450_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179963.4]
  reg [31:0] _RAND_394;
  reg  _T_451_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179966.4]
  reg [31:0] _RAND_395;
  reg  _T_452_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179969.4]
  reg [31:0] _RAND_396;
  reg  _T_453_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179972.4]
  reg [31:0] _RAND_397;
  reg  _T_454_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179975.4]
  reg [31:0] _RAND_398;
  reg  _T_455_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179978.4]
  reg [31:0] _RAND_399;
  reg  _T_456_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179981.4]
  reg [31:0] _RAND_400;
  reg  _T_457_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179984.4]
  reg [31:0] _RAND_401;
  reg  _T_458_0; // @[Mesh.scala 76:30:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179987.4]
  reg [31:0] _RAND_402;
  reg  _T_459_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179989.4]
  reg [31:0] _RAND_403;
  reg  _T_460_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179992.4]
  reg [31:0] _RAND_404;
  reg  _T_461_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179995.4]
  reg [31:0] _RAND_405;
  reg  _T_462_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179998.4]
  reg [31:0] _RAND_406;
  reg  _T_463_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180001.4]
  reg [31:0] _RAND_407;
  reg  _T_464_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180004.4]
  reg [31:0] _RAND_408;
  reg  _T_465_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180007.4]
  reg [31:0] _RAND_409;
  reg  _T_466_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180010.4]
  reg [31:0] _RAND_410;
  reg  _T_467_0; // @[Mesh.scala 76:30:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180013.4]
  reg [31:0] _RAND_411;
  reg  _T_468_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180015.4]
  reg [31:0] _RAND_412;
  reg  _T_469_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180018.4]
  reg [31:0] _RAND_413;
  reg  _T_470_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180021.4]
  reg [31:0] _RAND_414;
  reg  _T_471_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180024.4]
  reg [31:0] _RAND_415;
  reg  _T_472_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180027.4]
  reg [31:0] _RAND_416;
  reg  _T_473_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180030.4]
  reg [31:0] _RAND_417;
  reg  _T_474_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180033.4]
  reg [31:0] _RAND_418;
  reg  _T_475_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180036.4]
  reg [31:0] _RAND_419;
  reg  _T_476_0; // @[Mesh.scala 76:30:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180039.4]
  reg [31:0] _RAND_420;
  reg  _T_477_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180041.4]
  reg [31:0] _RAND_421;
  reg  _T_478_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180044.4]
  reg [31:0] _RAND_422;
  reg  _T_479_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180047.4]
  reg [31:0] _RAND_423;
  reg  _T_480_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180050.4]
  reg [31:0] _RAND_424;
  reg  _T_481_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180053.4]
  reg [31:0] _RAND_425;
  reg  _T_482_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180056.4]
  reg [31:0] _RAND_426;
  reg  _T_483_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180059.4]
  reg [31:0] _RAND_427;
  reg  _T_484_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180062.4]
  reg [31:0] _RAND_428;
  reg  _T_485_0; // @[Mesh.scala 76:30:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180065.4]
  reg [31:0] _RAND_429;
  reg  _T_486_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180067.4]
  reg [31:0] _RAND_430;
  reg  _T_487_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180070.4]
  reg [31:0] _RAND_431;
  reg  _T_488_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180073.4]
  reg [31:0] _RAND_432;
  reg  _T_489_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180076.4]
  reg [31:0] _RAND_433;
  reg  _T_490_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180079.4]
  reg [31:0] _RAND_434;
  reg  _T_491_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180082.4]
  reg [31:0] _RAND_435;
  reg  _T_492_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180085.4]
  reg [31:0] _RAND_436;
  reg  _T_493_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180088.4]
  reg [31:0] _RAND_437;
  reg  _T_494_0; // @[Mesh.scala 76:30:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180091.4]
  reg [31:0] _RAND_438;
  reg  _T_495_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180093.4]
  reg [31:0] _RAND_439;
  reg  _T_496_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180096.4]
  reg [31:0] _RAND_440;
  reg  _T_497_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180099.4]
  reg [31:0] _RAND_441;
  reg  _T_498_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180102.4]
  reg [31:0] _RAND_442;
  reg  _T_499_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180105.4]
  reg [31:0] _RAND_443;
  reg  _T_500_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180108.4]
  reg [31:0] _RAND_444;
  reg  _T_501_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180111.4]
  reg [31:0] _RAND_445;
  reg  _T_502_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180114.4]
  reg [31:0] _RAND_446;
  reg  _T_503_0; // @[Mesh.scala 76:30:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180117.4]
  reg [31:0] _RAND_447;
  reg  _T_504_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180119.4]
  reg [31:0] _RAND_448;
  reg  _T_505_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180122.4]
  reg [31:0] _RAND_449;
  reg  _T_506_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180125.4]
  reg [31:0] _RAND_450;
  reg  _T_507_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180128.4]
  reg [31:0] _RAND_451;
  reg  _T_508_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180131.4]
  reg [31:0] _RAND_452;
  reg  _T_509_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180134.4]
  reg [31:0] _RAND_453;
  reg  _T_510_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180137.4]
  reg [31:0] _RAND_454;
  reg  _T_511_0; // @[Mesh.scala 78:36:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180140.4]
  reg [31:0] _RAND_455;
  Tile mesh_0_0 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177823.4]
    .clock(mesh_0_0_clock),
    .io_in_a_0(mesh_0_0_io_in_a_0),
    .io_in_b_0(mesh_0_0_io_in_b_0),
    .io_in_d_0({`P_W'd0,{45{mesh_0_0_io_in_d_0[18]}},mesh_0_0_io_in_d_0}),
    .io_in_control_0_propagate(mesh_0_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_0_io_in_control_0_shift),
    .io_out_a_0(mesh_0_0_io_out_a_0),
    .io_out_c_0(mesh_0_0_io_out_c_0),
    .io_out_b_0(mesh_0_0_io_out_b_0),
    .io_out_control_0_propagate(mesh_0_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_0_io_out_control_0_shift),
    .io_in_valid_0(mesh_0_0_io_in_valid_0),
    .io_out_valid_0(mesh_0_0_io_out_valid_0)
  );
  Tile mesh_0_1 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177826.4]
    .clock(mesh_0_1_clock),
    .io_in_a_0(mesh_0_1_io_in_a_0),
    .io_in_b_0(mesh_0_1_io_in_b_0),
    .io_in_d_0({`P_W'd0,{45{mesh_0_1_io_in_d_0[18]}},mesh_0_1_io_in_d_0}),
    .io_in_control_0_propagate(mesh_0_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_1_io_in_control_0_shift),
    .io_out_a_0(mesh_0_1_io_out_a_0),
    .io_out_c_0(mesh_0_1_io_out_c_0),
    .io_out_b_0(mesh_0_1_io_out_b_0),
    .io_out_control_0_propagate(mesh_0_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_1_io_out_control_0_shift),
    .io_in_valid_0(mesh_0_1_io_in_valid_0),
    .io_out_valid_0(mesh_0_1_io_out_valid_0)
  );
  Tile mesh_0_2 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177829.4]
    .clock(mesh_0_2_clock),
    .io_in_a_0(mesh_0_2_io_in_a_0),
    .io_in_b_0(mesh_0_2_io_in_b_0),
    .io_in_d_0({`P_W'd0,{45{mesh_0_2_io_in_d_0[18]}},mesh_0_2_io_in_d_0}),
    .io_in_control_0_propagate(mesh_0_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_2_io_in_control_0_shift),
    .io_out_a_0(mesh_0_2_io_out_a_0),
    .io_out_c_0(mesh_0_2_io_out_c_0),
    .io_out_b_0(mesh_0_2_io_out_b_0),
    .io_out_control_0_propagate(mesh_0_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_2_io_out_control_0_shift),
    .io_in_valid_0(mesh_0_2_io_in_valid_0),
    .io_out_valid_0(mesh_0_2_io_out_valid_0)
  );
  Tile mesh_0_3 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177832.4]
    .clock(mesh_0_3_clock),
    .io_in_a_0(mesh_0_3_io_in_a_0),
    .io_in_b_0(mesh_0_3_io_in_b_0),
    .io_in_d_0({`P_W'd0,{45{mesh_0_3_io_in_d_0[18]}},mesh_0_3_io_in_d_0}),
    .io_in_control_0_propagate(mesh_0_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_3_io_in_control_0_shift),
    .io_out_a_0(mesh_0_3_io_out_a_0),
    .io_out_c_0(mesh_0_3_io_out_c_0),
    .io_out_b_0(mesh_0_3_io_out_b_0),
    .io_out_control_0_propagate(mesh_0_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_3_io_out_control_0_shift),
    .io_in_valid_0(mesh_0_3_io_in_valid_0),
    .io_out_valid_0(mesh_0_3_io_out_valid_0)
  );
  Tile mesh_0_4 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177835.4]
    .clock(mesh_0_4_clock),
    .io_in_a_0(mesh_0_4_io_in_a_0),
    .io_in_b_0(mesh_0_4_io_in_b_0),
    .io_in_d_0({`P_W'd0,{45{mesh_0_4_io_in_d_0[18]}},mesh_0_4_io_in_d_0}),
    .io_in_control_0_propagate(mesh_0_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_4_io_in_control_0_shift),
    .io_out_a_0(mesh_0_4_io_out_a_0),
    .io_out_c_0(mesh_0_4_io_out_c_0),
    .io_out_b_0(mesh_0_4_io_out_b_0),
    .io_out_control_0_propagate(mesh_0_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_4_io_out_control_0_shift),
    .io_in_valid_0(mesh_0_4_io_in_valid_0),
    .io_out_valid_0(mesh_0_4_io_out_valid_0)
  );
  Tile mesh_0_5 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177838.4]
    .clock(mesh_0_5_clock),
    .io_in_a_0(mesh_0_5_io_in_a_0),
    .io_in_b_0(mesh_0_5_io_in_b_0),
    .io_in_d_0({`P_W'd0,{45{mesh_0_5_io_in_d_0[18]}},mesh_0_5_io_in_d_0}),
    .io_in_control_0_propagate(mesh_0_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_5_io_in_control_0_shift),
    .io_out_a_0(mesh_0_5_io_out_a_0),
    .io_out_c_0(mesh_0_5_io_out_c_0),
    .io_out_b_0(mesh_0_5_io_out_b_0),
    .io_out_control_0_propagate(mesh_0_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_5_io_out_control_0_shift),
    .io_in_valid_0(mesh_0_5_io_in_valid_0),
    .io_out_valid_0(mesh_0_5_io_out_valid_0)
  );
  Tile mesh_0_6 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177841.4]
    .clock(mesh_0_6_clock),
    .io_in_a_0(mesh_0_6_io_in_a_0),
    .io_in_b_0(mesh_0_6_io_in_b_0),
    .io_in_d_0({`P_W'd0,{45{mesh_0_6_io_in_d_0[18]}},mesh_0_6_io_in_d_0}),
    .io_in_control_0_propagate(mesh_0_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_6_io_in_control_0_shift),
    .io_out_a_0(mesh_0_6_io_out_a_0),
    .io_out_c_0(mesh_0_6_io_out_c_0),
    .io_out_b_0(mesh_0_6_io_out_b_0),
    .io_out_control_0_propagate(mesh_0_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_6_io_out_control_0_shift),
    .io_in_valid_0(mesh_0_6_io_in_valid_0),
    .io_out_valid_0(mesh_0_6_io_out_valid_0)
  );
  Tile mesh_0_7 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177844.4]
    .clock(mesh_0_7_clock),
    .io_in_a_0(mesh_0_7_io_in_a_0),
    .io_in_b_0(mesh_0_7_io_in_b_0),
    .io_in_d_0({`P_W'd0,{45{mesh_0_7_io_in_d_0[18]}},mesh_0_7_io_in_d_0}),
    .io_in_control_0_propagate(mesh_0_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_0_7_io_in_control_0_shift),
    .io_out_a_0(mesh_0_7_io_out_a_0),
    .io_out_c_0(mesh_0_7_io_out_c_0),
    .io_out_b_0(mesh_0_7_io_out_b_0),
    .io_out_control_0_propagate(mesh_0_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_0_7_io_out_control_0_shift),
    .io_in_valid_0(mesh_0_7_io_in_valid_0),
    .io_out_valid_0(mesh_0_7_io_out_valid_0)
  );
  Tile mesh_1_0 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177847.4]
    .clock(mesh_1_0_clock),
    .io_in_a_0(mesh_1_0_io_in_a_0),
    .io_in_b_0(mesh_1_0_io_in_b_0),
    .io_in_d_0(mesh_1_0_io_in_d_0),
    .io_in_control_0_propagate(mesh_1_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_0_io_in_control_0_shift),
    .io_out_a_0(mesh_1_0_io_out_a_0),
    .io_out_c_0(mesh_1_0_io_out_c_0),
    .io_out_b_0(mesh_1_0_io_out_b_0),
    .io_out_control_0_propagate(mesh_1_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_0_io_out_control_0_shift),
    .io_in_valid_0(mesh_1_0_io_in_valid_0),
    .io_out_valid_0(mesh_1_0_io_out_valid_0)
  );
  Tile mesh_1_1 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177850.4]
    .clock(mesh_1_1_clock),
    .io_in_a_0(mesh_1_1_io_in_a_0),
    .io_in_b_0(mesh_1_1_io_in_b_0),
    .io_in_d_0(mesh_1_1_io_in_d_0),
    .io_in_control_0_propagate(mesh_1_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_1_io_in_control_0_shift),
    .io_out_a_0(mesh_1_1_io_out_a_0),
    .io_out_c_0(mesh_1_1_io_out_c_0),
    .io_out_b_0(mesh_1_1_io_out_b_0),
    .io_out_control_0_propagate(mesh_1_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_1_io_out_control_0_shift),
    .io_in_valid_0(mesh_1_1_io_in_valid_0),
    .io_out_valid_0(mesh_1_1_io_out_valid_0)
  );
  Tile mesh_1_2 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177853.4]
    .clock(mesh_1_2_clock),
    .io_in_a_0(mesh_1_2_io_in_a_0),
    .io_in_b_0(mesh_1_2_io_in_b_0),
    .io_in_d_0(mesh_1_2_io_in_d_0),
    .io_in_control_0_propagate(mesh_1_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_2_io_in_control_0_shift),
    .io_out_a_0(mesh_1_2_io_out_a_0),
    .io_out_c_0(mesh_1_2_io_out_c_0),
    .io_out_b_0(mesh_1_2_io_out_b_0),
    .io_out_control_0_propagate(mesh_1_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_2_io_out_control_0_shift),
    .io_in_valid_0(mesh_1_2_io_in_valid_0),
    .io_out_valid_0(mesh_1_2_io_out_valid_0)
  );
  Tile mesh_1_3 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177856.4]
    .clock(mesh_1_3_clock),
    .io_in_a_0(mesh_1_3_io_in_a_0),
    .io_in_b_0(mesh_1_3_io_in_b_0),
    .io_in_d_0(mesh_1_3_io_in_d_0),
    .io_in_control_0_propagate(mesh_1_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_3_io_in_control_0_shift),
    .io_out_a_0(mesh_1_3_io_out_a_0),
    .io_out_c_0(mesh_1_3_io_out_c_0),
    .io_out_b_0(mesh_1_3_io_out_b_0),
    .io_out_control_0_propagate(mesh_1_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_3_io_out_control_0_shift),
    .io_in_valid_0(mesh_1_3_io_in_valid_0),
    .io_out_valid_0(mesh_1_3_io_out_valid_0)
  );
  Tile mesh_1_4 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177859.4]
    .clock(mesh_1_4_clock),
    .io_in_a_0(mesh_1_4_io_in_a_0),
    .io_in_b_0(mesh_1_4_io_in_b_0),
    .io_in_d_0(mesh_1_4_io_in_d_0),
    .io_in_control_0_propagate(mesh_1_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_4_io_in_control_0_shift),
    .io_out_a_0(mesh_1_4_io_out_a_0),
    .io_out_c_0(mesh_1_4_io_out_c_0),
    .io_out_b_0(mesh_1_4_io_out_b_0),
    .io_out_control_0_propagate(mesh_1_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_4_io_out_control_0_shift),
    .io_in_valid_0(mesh_1_4_io_in_valid_0),
    .io_out_valid_0(mesh_1_4_io_out_valid_0)
  );
  Tile mesh_1_5 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177862.4]
    .clock(mesh_1_5_clock),
    .io_in_a_0(mesh_1_5_io_in_a_0),
    .io_in_b_0(mesh_1_5_io_in_b_0),
    .io_in_d_0(mesh_1_5_io_in_d_0),
    .io_in_control_0_propagate(mesh_1_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_5_io_in_control_0_shift),
    .io_out_a_0(mesh_1_5_io_out_a_0),
    .io_out_c_0(mesh_1_5_io_out_c_0),
    .io_out_b_0(mesh_1_5_io_out_b_0),
    .io_out_control_0_propagate(mesh_1_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_5_io_out_control_0_shift),
    .io_in_valid_0(mesh_1_5_io_in_valid_0),
    .io_out_valid_0(mesh_1_5_io_out_valid_0)
  );
  Tile mesh_1_6 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177865.4]
    .clock(mesh_1_6_clock),
    .io_in_a_0(mesh_1_6_io_in_a_0),
    .io_in_b_0(mesh_1_6_io_in_b_0),
    .io_in_d_0(mesh_1_6_io_in_d_0),
    .io_in_control_0_propagate(mesh_1_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_6_io_in_control_0_shift),
    .io_out_a_0(mesh_1_6_io_out_a_0),
    .io_out_c_0(mesh_1_6_io_out_c_0),
    .io_out_b_0(mesh_1_6_io_out_b_0),
    .io_out_control_0_propagate(mesh_1_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_6_io_out_control_0_shift),
    .io_in_valid_0(mesh_1_6_io_in_valid_0),
    .io_out_valid_0(mesh_1_6_io_out_valid_0)
  );
  Tile mesh_1_7 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177868.4]
    .clock(mesh_1_7_clock),
    .io_in_a_0(mesh_1_7_io_in_a_0),
    .io_in_b_0(mesh_1_7_io_in_b_0),
    .io_in_d_0(mesh_1_7_io_in_d_0),
    .io_in_control_0_propagate(mesh_1_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_1_7_io_in_control_0_shift),
    .io_out_a_0(mesh_1_7_io_out_a_0),
    .io_out_c_0(mesh_1_7_io_out_c_0),
    .io_out_b_0(mesh_1_7_io_out_b_0),
    .io_out_control_0_propagate(mesh_1_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_1_7_io_out_control_0_shift),
    .io_in_valid_0(mesh_1_7_io_in_valid_0),
    .io_out_valid_0(mesh_1_7_io_out_valid_0)
  );
  Tile mesh_2_0 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177871.4]
    .clock(mesh_2_0_clock),
    .io_in_a_0(mesh_2_0_io_in_a_0),
    .io_in_b_0(mesh_2_0_io_in_b_0),
    .io_in_d_0(mesh_2_0_io_in_d_0),
    .io_in_control_0_propagate(mesh_2_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_0_io_in_control_0_shift),
    .io_out_a_0(mesh_2_0_io_out_a_0),
    .io_out_c_0(mesh_2_0_io_out_c_0),
    .io_out_b_0(mesh_2_0_io_out_b_0),
    .io_out_control_0_propagate(mesh_2_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_0_io_out_control_0_shift),
    .io_in_valid_0(mesh_2_0_io_in_valid_0),
    .io_out_valid_0(mesh_2_0_io_out_valid_0)
  );
  Tile mesh_2_1 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177874.4]
    .clock(mesh_2_1_clock),
    .io_in_a_0(mesh_2_1_io_in_a_0),
    .io_in_b_0(mesh_2_1_io_in_b_0),
    .io_in_d_0(mesh_2_1_io_in_d_0),
    .io_in_control_0_propagate(mesh_2_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_1_io_in_control_0_shift),
    .io_out_a_0(mesh_2_1_io_out_a_0),
    .io_out_c_0(mesh_2_1_io_out_c_0),
    .io_out_b_0(mesh_2_1_io_out_b_0),
    .io_out_control_0_propagate(mesh_2_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_1_io_out_control_0_shift),
    .io_in_valid_0(mesh_2_1_io_in_valid_0),
    .io_out_valid_0(mesh_2_1_io_out_valid_0)
  );
  Tile mesh_2_2 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177877.4]
    .clock(mesh_2_2_clock),
    .io_in_a_0(mesh_2_2_io_in_a_0),
    .io_in_b_0(mesh_2_2_io_in_b_0),
    .io_in_d_0(mesh_2_2_io_in_d_0),
    .io_in_control_0_propagate(mesh_2_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_2_io_in_control_0_shift),
    .io_out_a_0(mesh_2_2_io_out_a_0),
    .io_out_c_0(mesh_2_2_io_out_c_0),
    .io_out_b_0(mesh_2_2_io_out_b_0),
    .io_out_control_0_propagate(mesh_2_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_2_io_out_control_0_shift),
    .io_in_valid_0(mesh_2_2_io_in_valid_0),
    .io_out_valid_0(mesh_2_2_io_out_valid_0)
  );
  Tile mesh_2_3 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177880.4]
    .clock(mesh_2_3_clock),
    .io_in_a_0(mesh_2_3_io_in_a_0),
    .io_in_b_0(mesh_2_3_io_in_b_0),
    .io_in_d_0(mesh_2_3_io_in_d_0),
    .io_in_control_0_propagate(mesh_2_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_3_io_in_control_0_shift),
    .io_out_a_0(mesh_2_3_io_out_a_0),
    .io_out_c_0(mesh_2_3_io_out_c_0),
    .io_out_b_0(mesh_2_3_io_out_b_0),
    .io_out_control_0_propagate(mesh_2_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_3_io_out_control_0_shift),
    .io_in_valid_0(mesh_2_3_io_in_valid_0),
    .io_out_valid_0(mesh_2_3_io_out_valid_0)
  );
  Tile mesh_2_4 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177883.4]
    .clock(mesh_2_4_clock),
    .io_in_a_0(mesh_2_4_io_in_a_0),
    .io_in_b_0(mesh_2_4_io_in_b_0),
    .io_in_d_0(mesh_2_4_io_in_d_0),
    .io_in_control_0_propagate(mesh_2_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_4_io_in_control_0_shift),
    .io_out_a_0(mesh_2_4_io_out_a_0),
    .io_out_c_0(mesh_2_4_io_out_c_0),
    .io_out_b_0(mesh_2_4_io_out_b_0),
    .io_out_control_0_propagate(mesh_2_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_4_io_out_control_0_shift),
    .io_in_valid_0(mesh_2_4_io_in_valid_0),
    .io_out_valid_0(mesh_2_4_io_out_valid_0)
  );
  Tile mesh_2_5 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177886.4]
    .clock(mesh_2_5_clock),
    .io_in_a_0(mesh_2_5_io_in_a_0),
    .io_in_b_0(mesh_2_5_io_in_b_0),
    .io_in_d_0(mesh_2_5_io_in_d_0),
    .io_in_control_0_propagate(mesh_2_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_5_io_in_control_0_shift),
    .io_out_a_0(mesh_2_5_io_out_a_0),
    .io_out_c_0(mesh_2_5_io_out_c_0),
    .io_out_b_0(mesh_2_5_io_out_b_0),
    .io_out_control_0_propagate(mesh_2_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_5_io_out_control_0_shift),
    .io_in_valid_0(mesh_2_5_io_in_valid_0),
    .io_out_valid_0(mesh_2_5_io_out_valid_0)
  );
  Tile mesh_2_6 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177889.4]
    .clock(mesh_2_6_clock),
    .io_in_a_0(mesh_2_6_io_in_a_0),
    .io_in_b_0(mesh_2_6_io_in_b_0),
    .io_in_d_0(mesh_2_6_io_in_d_0),
    .io_in_control_0_propagate(mesh_2_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_6_io_in_control_0_shift),
    .io_out_a_0(mesh_2_6_io_out_a_0),
    .io_out_c_0(mesh_2_6_io_out_c_0),
    .io_out_b_0(mesh_2_6_io_out_b_0),
    .io_out_control_0_propagate(mesh_2_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_6_io_out_control_0_shift),
    .io_in_valid_0(mesh_2_6_io_in_valid_0),
    .io_out_valid_0(mesh_2_6_io_out_valid_0)
  );
  Tile mesh_2_7 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177892.4]
    .clock(mesh_2_7_clock),
    .io_in_a_0(mesh_2_7_io_in_a_0),
    .io_in_b_0(mesh_2_7_io_in_b_0),
    .io_in_d_0(mesh_2_7_io_in_d_0),
    .io_in_control_0_propagate(mesh_2_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_2_7_io_in_control_0_shift),
    .io_out_a_0(mesh_2_7_io_out_a_0),
    .io_out_c_0(mesh_2_7_io_out_c_0),
    .io_out_b_0(mesh_2_7_io_out_b_0),
    .io_out_control_0_propagate(mesh_2_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_2_7_io_out_control_0_shift),
    .io_in_valid_0(mesh_2_7_io_in_valid_0),
    .io_out_valid_0(mesh_2_7_io_out_valid_0)
  );
  Tile mesh_3_0 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177895.4]
    .clock(mesh_3_0_clock),
    .io_in_a_0(mesh_3_0_io_in_a_0),
    .io_in_b_0(mesh_3_0_io_in_b_0),
    .io_in_d_0(mesh_3_0_io_in_d_0),
    .io_in_control_0_propagate(mesh_3_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_0_io_in_control_0_shift),
    .io_out_a_0(mesh_3_0_io_out_a_0),
    .io_out_c_0(mesh_3_0_io_out_c_0),
    .io_out_b_0(mesh_3_0_io_out_b_0),
    .io_out_control_0_propagate(mesh_3_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_0_io_out_control_0_shift),
    .io_in_valid_0(mesh_3_0_io_in_valid_0),
    .io_out_valid_0(mesh_3_0_io_out_valid_0)
  );
  Tile mesh_3_1 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177898.4]
    .clock(mesh_3_1_clock),
    .io_in_a_0(mesh_3_1_io_in_a_0),
    .io_in_b_0(mesh_3_1_io_in_b_0),
    .io_in_d_0(mesh_3_1_io_in_d_0),
    .io_in_control_0_propagate(mesh_3_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_1_io_in_control_0_shift),
    .io_out_a_0(mesh_3_1_io_out_a_0),
    .io_out_c_0(mesh_3_1_io_out_c_0),
    .io_out_b_0(mesh_3_1_io_out_b_0),
    .io_out_control_0_propagate(mesh_3_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_1_io_out_control_0_shift),
    .io_in_valid_0(mesh_3_1_io_in_valid_0),
    .io_out_valid_0(mesh_3_1_io_out_valid_0)
  );
  Tile mesh_3_2 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177901.4]
    .clock(mesh_3_2_clock),
    .io_in_a_0(mesh_3_2_io_in_a_0),
    .io_in_b_0(mesh_3_2_io_in_b_0),
    .io_in_d_0(mesh_3_2_io_in_d_0),
    .io_in_control_0_propagate(mesh_3_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_2_io_in_control_0_shift),
    .io_out_a_0(mesh_3_2_io_out_a_0),
    .io_out_c_0(mesh_3_2_io_out_c_0),
    .io_out_b_0(mesh_3_2_io_out_b_0),
    .io_out_control_0_propagate(mesh_3_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_2_io_out_control_0_shift),
    .io_in_valid_0(mesh_3_2_io_in_valid_0),
    .io_out_valid_0(mesh_3_2_io_out_valid_0)
  );
  Tile mesh_3_3 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177904.4]
    .clock(mesh_3_3_clock),
    .io_in_a_0(mesh_3_3_io_in_a_0),
    .io_in_b_0(mesh_3_3_io_in_b_0),
    .io_in_d_0(mesh_3_3_io_in_d_0),
    .io_in_control_0_propagate(mesh_3_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_3_io_in_control_0_shift),
    .io_out_a_0(mesh_3_3_io_out_a_0),
    .io_out_c_0(mesh_3_3_io_out_c_0),
    .io_out_b_0(mesh_3_3_io_out_b_0),
    .io_out_control_0_propagate(mesh_3_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_3_io_out_control_0_shift),
    .io_in_valid_0(mesh_3_3_io_in_valid_0),
    .io_out_valid_0(mesh_3_3_io_out_valid_0)
  );
  Tile mesh_3_4 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177907.4]
    .clock(mesh_3_4_clock),
    .io_in_a_0(mesh_3_4_io_in_a_0),
    .io_in_b_0(mesh_3_4_io_in_b_0),
    .io_in_d_0(mesh_3_4_io_in_d_0),
    .io_in_control_0_propagate(mesh_3_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_4_io_in_control_0_shift),
    .io_out_a_0(mesh_3_4_io_out_a_0),
    .io_out_c_0(mesh_3_4_io_out_c_0),
    .io_out_b_0(mesh_3_4_io_out_b_0),
    .io_out_control_0_propagate(mesh_3_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_4_io_out_control_0_shift),
    .io_in_valid_0(mesh_3_4_io_in_valid_0),
    .io_out_valid_0(mesh_3_4_io_out_valid_0)
  );
  Tile mesh_3_5 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177910.4]
    .clock(mesh_3_5_clock),
    .io_in_a_0(mesh_3_5_io_in_a_0),
    .io_in_b_0(mesh_3_5_io_in_b_0),
    .io_in_d_0(mesh_3_5_io_in_d_0),
    .io_in_control_0_propagate(mesh_3_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_5_io_in_control_0_shift),
    .io_out_a_0(mesh_3_5_io_out_a_0),
    .io_out_c_0(mesh_3_5_io_out_c_0),
    .io_out_b_0(mesh_3_5_io_out_b_0),
    .io_out_control_0_propagate(mesh_3_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_5_io_out_control_0_shift),
    .io_in_valid_0(mesh_3_5_io_in_valid_0),
    .io_out_valid_0(mesh_3_5_io_out_valid_0)
  );
  Tile mesh_3_6 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177913.4]
    .clock(mesh_3_6_clock),
    .io_in_a_0(mesh_3_6_io_in_a_0),
    .io_in_b_0(mesh_3_6_io_in_b_0),
    .io_in_d_0(mesh_3_6_io_in_d_0),
    .io_in_control_0_propagate(mesh_3_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_6_io_in_control_0_shift),
    .io_out_a_0(mesh_3_6_io_out_a_0),
    .io_out_c_0(mesh_3_6_io_out_c_0),
    .io_out_b_0(mesh_3_6_io_out_b_0),
    .io_out_control_0_propagate(mesh_3_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_6_io_out_control_0_shift),
    .io_in_valid_0(mesh_3_6_io_in_valid_0),
    .io_out_valid_0(mesh_3_6_io_out_valid_0)
  );
  Tile mesh_3_7 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177916.4]
    .clock(mesh_3_7_clock),
    .io_in_a_0(mesh_3_7_io_in_a_0),
    .io_in_b_0(mesh_3_7_io_in_b_0),
    .io_in_d_0(mesh_3_7_io_in_d_0),
    .io_in_control_0_propagate(mesh_3_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_3_7_io_in_control_0_shift),
    .io_out_a_0(mesh_3_7_io_out_a_0),
    .io_out_c_0(mesh_3_7_io_out_c_0),
    .io_out_b_0(mesh_3_7_io_out_b_0),
    .io_out_control_0_propagate(mesh_3_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_3_7_io_out_control_0_shift),
    .io_in_valid_0(mesh_3_7_io_in_valid_0),
    .io_out_valid_0(mesh_3_7_io_out_valid_0)
  );
  Tile mesh_4_0 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177919.4]
    .clock(mesh_4_0_clock),
    .io_in_a_0(mesh_4_0_io_in_a_0),
    .io_in_b_0(mesh_4_0_io_in_b_0),
    .io_in_d_0(mesh_4_0_io_in_d_0),
    .io_in_control_0_propagate(mesh_4_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_0_io_in_control_0_shift),
    .io_out_a_0(mesh_4_0_io_out_a_0),
    .io_out_c_0(mesh_4_0_io_out_c_0),
    .io_out_b_0(mesh_4_0_io_out_b_0),
    .io_out_control_0_propagate(mesh_4_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_0_io_out_control_0_shift),
    .io_in_valid_0(mesh_4_0_io_in_valid_0),
    .io_out_valid_0(mesh_4_0_io_out_valid_0)
  );
  Tile mesh_4_1 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177922.4]
    .clock(mesh_4_1_clock),
    .io_in_a_0(mesh_4_1_io_in_a_0),
    .io_in_b_0(mesh_4_1_io_in_b_0),
    .io_in_d_0(mesh_4_1_io_in_d_0),
    .io_in_control_0_propagate(mesh_4_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_1_io_in_control_0_shift),
    .io_out_a_0(mesh_4_1_io_out_a_0),
    .io_out_c_0(mesh_4_1_io_out_c_0),
    .io_out_b_0(mesh_4_1_io_out_b_0),
    .io_out_control_0_propagate(mesh_4_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_1_io_out_control_0_shift),
    .io_in_valid_0(mesh_4_1_io_in_valid_0),
    .io_out_valid_0(mesh_4_1_io_out_valid_0)
  );
  Tile mesh_4_2 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177925.4]
    .clock(mesh_4_2_clock),
    .io_in_a_0(mesh_4_2_io_in_a_0),
    .io_in_b_0(mesh_4_2_io_in_b_0),
    .io_in_d_0(mesh_4_2_io_in_d_0),
    .io_in_control_0_propagate(mesh_4_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_2_io_in_control_0_shift),
    .io_out_a_0(mesh_4_2_io_out_a_0),
    .io_out_c_0(mesh_4_2_io_out_c_0),
    .io_out_b_0(mesh_4_2_io_out_b_0),
    .io_out_control_0_propagate(mesh_4_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_2_io_out_control_0_shift),
    .io_in_valid_0(mesh_4_2_io_in_valid_0),
    .io_out_valid_0(mesh_4_2_io_out_valid_0)
  );
  Tile mesh_4_3 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177928.4]
    .clock(mesh_4_3_clock),
    .io_in_a_0(mesh_4_3_io_in_a_0),
    .io_in_b_0(mesh_4_3_io_in_b_0),
    .io_in_d_0(mesh_4_3_io_in_d_0),
    .io_in_control_0_propagate(mesh_4_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_3_io_in_control_0_shift),
    .io_out_a_0(mesh_4_3_io_out_a_0),
    .io_out_c_0(mesh_4_3_io_out_c_0),
    .io_out_b_0(mesh_4_3_io_out_b_0),
    .io_out_control_0_propagate(mesh_4_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_3_io_out_control_0_shift),
    .io_in_valid_0(mesh_4_3_io_in_valid_0),
    .io_out_valid_0(mesh_4_3_io_out_valid_0)
  );
  Tile mesh_4_4 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177931.4]
    .clock(mesh_4_4_clock),
    .io_in_a_0(mesh_4_4_io_in_a_0),
    .io_in_b_0(mesh_4_4_io_in_b_0),
    .io_in_d_0(mesh_4_4_io_in_d_0),
    .io_in_control_0_propagate(mesh_4_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_4_io_in_control_0_shift),
    .io_out_a_0(mesh_4_4_io_out_a_0),
    .io_out_c_0(mesh_4_4_io_out_c_0),
    .io_out_b_0(mesh_4_4_io_out_b_0),
    .io_out_control_0_propagate(mesh_4_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_4_io_out_control_0_shift),
    .io_in_valid_0(mesh_4_4_io_in_valid_0),
    .io_out_valid_0(mesh_4_4_io_out_valid_0)
  );
  Tile mesh_4_5 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177934.4]
    .clock(mesh_4_5_clock),
    .io_in_a_0(mesh_4_5_io_in_a_0),
    .io_in_b_0(mesh_4_5_io_in_b_0),
    .io_in_d_0(mesh_4_5_io_in_d_0),
    .io_in_control_0_propagate(mesh_4_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_5_io_in_control_0_shift),
    .io_out_a_0(mesh_4_5_io_out_a_0),
    .io_out_c_0(mesh_4_5_io_out_c_0),
    .io_out_b_0(mesh_4_5_io_out_b_0),
    .io_out_control_0_propagate(mesh_4_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_5_io_out_control_0_shift),
    .io_in_valid_0(mesh_4_5_io_in_valid_0),
    .io_out_valid_0(mesh_4_5_io_out_valid_0)
  );
  Tile mesh_4_6 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177937.4]
    .clock(mesh_4_6_clock),
    .io_in_a_0(mesh_4_6_io_in_a_0),
    .io_in_b_0(mesh_4_6_io_in_b_0),
    .io_in_d_0(mesh_4_6_io_in_d_0),
    .io_in_control_0_propagate(mesh_4_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_6_io_in_control_0_shift),
    .io_out_a_0(mesh_4_6_io_out_a_0),
    .io_out_c_0(mesh_4_6_io_out_c_0),
    .io_out_b_0(mesh_4_6_io_out_b_0),
    .io_out_control_0_propagate(mesh_4_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_6_io_out_control_0_shift),
    .io_in_valid_0(mesh_4_6_io_in_valid_0),
    .io_out_valid_0(mesh_4_6_io_out_valid_0)
  );
  Tile mesh_4_7 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177940.4]
    .clock(mesh_4_7_clock),
    .io_in_a_0(mesh_4_7_io_in_a_0),
    .io_in_b_0(mesh_4_7_io_in_b_0),
    .io_in_d_0(mesh_4_7_io_in_d_0),
    .io_in_control_0_propagate(mesh_4_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_4_7_io_in_control_0_shift),
    .io_out_a_0(mesh_4_7_io_out_a_0),
    .io_out_c_0(mesh_4_7_io_out_c_0),
    .io_out_b_0(mesh_4_7_io_out_b_0),
    .io_out_control_0_propagate(mesh_4_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_4_7_io_out_control_0_shift),
    .io_in_valid_0(mesh_4_7_io_in_valid_0),
    .io_out_valid_0(mesh_4_7_io_out_valid_0)
  );
  Tile mesh_5_0 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177943.4]
    .clock(mesh_5_0_clock),
    .io_in_a_0(mesh_5_0_io_in_a_0),
    .io_in_b_0(mesh_5_0_io_in_b_0),
    .io_in_d_0(mesh_5_0_io_in_d_0),
    .io_in_control_0_propagate(mesh_5_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_0_io_in_control_0_shift),
    .io_out_a_0(mesh_5_0_io_out_a_0),
    .io_out_c_0(mesh_5_0_io_out_c_0),
    .io_out_b_0(mesh_5_0_io_out_b_0),
    .io_out_control_0_propagate(mesh_5_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_0_io_out_control_0_shift),
    .io_in_valid_0(mesh_5_0_io_in_valid_0),
    .io_out_valid_0(mesh_5_0_io_out_valid_0)
  );
  Tile mesh_5_1 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177946.4]
    .clock(mesh_5_1_clock),
    .io_in_a_0(mesh_5_1_io_in_a_0),
    .io_in_b_0(mesh_5_1_io_in_b_0),
    .io_in_d_0(mesh_5_1_io_in_d_0),
    .io_in_control_0_propagate(mesh_5_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_1_io_in_control_0_shift),
    .io_out_a_0(mesh_5_1_io_out_a_0),
    .io_out_c_0(mesh_5_1_io_out_c_0),
    .io_out_b_0(mesh_5_1_io_out_b_0),
    .io_out_control_0_propagate(mesh_5_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_1_io_out_control_0_shift),
    .io_in_valid_0(mesh_5_1_io_in_valid_0),
    .io_out_valid_0(mesh_5_1_io_out_valid_0)
  );
  Tile mesh_5_2 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177949.4]
    .clock(mesh_5_2_clock),
    .io_in_a_0(mesh_5_2_io_in_a_0),
    .io_in_b_0(mesh_5_2_io_in_b_0),
    .io_in_d_0(mesh_5_2_io_in_d_0),
    .io_in_control_0_propagate(mesh_5_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_2_io_in_control_0_shift),
    .io_out_a_0(mesh_5_2_io_out_a_0),
    .io_out_c_0(mesh_5_2_io_out_c_0),
    .io_out_b_0(mesh_5_2_io_out_b_0),
    .io_out_control_0_propagate(mesh_5_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_2_io_out_control_0_shift),
    .io_in_valid_0(mesh_5_2_io_in_valid_0),
    .io_out_valid_0(mesh_5_2_io_out_valid_0)
  );
  Tile mesh_5_3 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177952.4]
    .clock(mesh_5_3_clock),
    .io_in_a_0(mesh_5_3_io_in_a_0),
    .io_in_b_0(mesh_5_3_io_in_b_0),
    .io_in_d_0(mesh_5_3_io_in_d_0),
    .io_in_control_0_propagate(mesh_5_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_3_io_in_control_0_shift),
    .io_out_a_0(mesh_5_3_io_out_a_0),
    .io_out_c_0(mesh_5_3_io_out_c_0),
    .io_out_b_0(mesh_5_3_io_out_b_0),
    .io_out_control_0_propagate(mesh_5_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_3_io_out_control_0_shift),
    .io_in_valid_0(mesh_5_3_io_in_valid_0),
    .io_out_valid_0(mesh_5_3_io_out_valid_0)
  );
  Tile mesh_5_4 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177955.4]
    .clock(mesh_5_4_clock),
    .io_in_a_0(mesh_5_4_io_in_a_0),
    .io_in_b_0(mesh_5_4_io_in_b_0),
    .io_in_d_0(mesh_5_4_io_in_d_0),
    .io_in_control_0_propagate(mesh_5_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_4_io_in_control_0_shift),
    .io_out_a_0(mesh_5_4_io_out_a_0),
    .io_out_c_0(mesh_5_4_io_out_c_0),
    .io_out_b_0(mesh_5_4_io_out_b_0),
    .io_out_control_0_propagate(mesh_5_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_4_io_out_control_0_shift),
    .io_in_valid_0(mesh_5_4_io_in_valid_0),
    .io_out_valid_0(mesh_5_4_io_out_valid_0)
  );
  Tile mesh_5_5 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177958.4]
    .clock(mesh_5_5_clock),
    .io_in_a_0(mesh_5_5_io_in_a_0),
    .io_in_b_0(mesh_5_5_io_in_b_0),
    .io_in_d_0(mesh_5_5_io_in_d_0),
    .io_in_control_0_propagate(mesh_5_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_5_io_in_control_0_shift),
    .io_out_a_0(mesh_5_5_io_out_a_0),
    .io_out_c_0(mesh_5_5_io_out_c_0),
    .io_out_b_0(mesh_5_5_io_out_b_0),
    .io_out_control_0_propagate(mesh_5_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_5_io_out_control_0_shift),
    .io_in_valid_0(mesh_5_5_io_in_valid_0),
    .io_out_valid_0(mesh_5_5_io_out_valid_0)
  );
  Tile mesh_5_6 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177961.4]
    .clock(mesh_5_6_clock),
    .io_in_a_0(mesh_5_6_io_in_a_0),
    .io_in_b_0(mesh_5_6_io_in_b_0),
    .io_in_d_0(mesh_5_6_io_in_d_0),
    .io_in_control_0_propagate(mesh_5_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_6_io_in_control_0_shift),
    .io_out_a_0(mesh_5_6_io_out_a_0),
    .io_out_c_0(mesh_5_6_io_out_c_0),
    .io_out_b_0(mesh_5_6_io_out_b_0),
    .io_out_control_0_propagate(mesh_5_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_6_io_out_control_0_shift),
    .io_in_valid_0(mesh_5_6_io_in_valid_0),
    .io_out_valid_0(mesh_5_6_io_out_valid_0)
  );
  Tile mesh_5_7 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177964.4]
    .clock(mesh_5_7_clock),
    .io_in_a_0(mesh_5_7_io_in_a_0),
    .io_in_b_0(mesh_5_7_io_in_b_0),
    .io_in_d_0(mesh_5_7_io_in_d_0),
    .io_in_control_0_propagate(mesh_5_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_5_7_io_in_control_0_shift),
    .io_out_a_0(mesh_5_7_io_out_a_0),
    .io_out_c_0(mesh_5_7_io_out_c_0),
    .io_out_b_0(mesh_5_7_io_out_b_0),
    .io_out_control_0_propagate(mesh_5_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_5_7_io_out_control_0_shift),
    .io_in_valid_0(mesh_5_7_io_in_valid_0),
    .io_out_valid_0(mesh_5_7_io_out_valid_0)
  );
  Tile mesh_6_0 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177967.4]
    .clock(mesh_6_0_clock),
    .io_in_a_0(mesh_6_0_io_in_a_0),
    .io_in_b_0(mesh_6_0_io_in_b_0),
    .io_in_d_0(mesh_6_0_io_in_d_0),
    .io_in_control_0_propagate(mesh_6_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_0_io_in_control_0_shift),
    .io_out_a_0(mesh_6_0_io_out_a_0),
    .io_out_c_0(mesh_6_0_io_out_c_0),
    .io_out_b_0(mesh_6_0_io_out_b_0),
    .io_out_control_0_propagate(mesh_6_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_0_io_out_control_0_shift),
    .io_in_valid_0(mesh_6_0_io_in_valid_0),
    .io_out_valid_0(mesh_6_0_io_out_valid_0)
  );
  Tile mesh_6_1 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177970.4]
    .clock(mesh_6_1_clock),
    .io_in_a_0(mesh_6_1_io_in_a_0),
    .io_in_b_0(mesh_6_1_io_in_b_0),
    .io_in_d_0(mesh_6_1_io_in_d_0),
    .io_in_control_0_propagate(mesh_6_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_1_io_in_control_0_shift),
    .io_out_a_0(mesh_6_1_io_out_a_0),
    .io_out_c_0(mesh_6_1_io_out_c_0),
    .io_out_b_0(mesh_6_1_io_out_b_0),
    .io_out_control_0_propagate(mesh_6_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_1_io_out_control_0_shift),
    .io_in_valid_0(mesh_6_1_io_in_valid_0),
    .io_out_valid_0(mesh_6_1_io_out_valid_0)
  );
  Tile mesh_6_2 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177973.4]
    .clock(mesh_6_2_clock),
    .io_in_a_0(mesh_6_2_io_in_a_0),
    .io_in_b_0(mesh_6_2_io_in_b_0),
    .io_in_d_0(mesh_6_2_io_in_d_0),
    .io_in_control_0_propagate(mesh_6_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_2_io_in_control_0_shift),
    .io_out_a_0(mesh_6_2_io_out_a_0),
    .io_out_c_0(mesh_6_2_io_out_c_0),
    .io_out_b_0(mesh_6_2_io_out_b_0),
    .io_out_control_0_propagate(mesh_6_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_2_io_out_control_0_shift),
    .io_in_valid_0(mesh_6_2_io_in_valid_0),
    .io_out_valid_0(mesh_6_2_io_out_valid_0)
  );
  Tile mesh_6_3 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177976.4]
    .clock(mesh_6_3_clock),
    .io_in_a_0(mesh_6_3_io_in_a_0),
    .io_in_b_0(mesh_6_3_io_in_b_0),
    .io_in_d_0(mesh_6_3_io_in_d_0),
    .io_in_control_0_propagate(mesh_6_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_3_io_in_control_0_shift),
    .io_out_a_0(mesh_6_3_io_out_a_0),
    .io_out_c_0(mesh_6_3_io_out_c_0),
    .io_out_b_0(mesh_6_3_io_out_b_0),
    .io_out_control_0_propagate(mesh_6_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_3_io_out_control_0_shift),
    .io_in_valid_0(mesh_6_3_io_in_valid_0),
    .io_out_valid_0(mesh_6_3_io_out_valid_0)
  );
  Tile mesh_6_4 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177979.4]
    .clock(mesh_6_4_clock),
    .io_in_a_0(mesh_6_4_io_in_a_0),
    .io_in_b_0(mesh_6_4_io_in_b_0),
    .io_in_d_0(mesh_6_4_io_in_d_0),
    .io_in_control_0_propagate(mesh_6_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_4_io_in_control_0_shift),
    .io_out_a_0(mesh_6_4_io_out_a_0),
    .io_out_c_0(mesh_6_4_io_out_c_0),
    .io_out_b_0(mesh_6_4_io_out_b_0),
    .io_out_control_0_propagate(mesh_6_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_4_io_out_control_0_shift),
    .io_in_valid_0(mesh_6_4_io_in_valid_0),
    .io_out_valid_0(mesh_6_4_io_out_valid_0)
  );
  Tile mesh_6_5 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177982.4]
    .clock(mesh_6_5_clock),
    .io_in_a_0(mesh_6_5_io_in_a_0),
    .io_in_b_0(mesh_6_5_io_in_b_0),
    .io_in_d_0(mesh_6_5_io_in_d_0),
    .io_in_control_0_propagate(mesh_6_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_5_io_in_control_0_shift),
    .io_out_a_0(mesh_6_5_io_out_a_0),
    .io_out_c_0(mesh_6_5_io_out_c_0),
    .io_out_b_0(mesh_6_5_io_out_b_0),
    .io_out_control_0_propagate(mesh_6_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_5_io_out_control_0_shift),
    .io_in_valid_0(mesh_6_5_io_in_valid_0),
    .io_out_valid_0(mesh_6_5_io_out_valid_0)
  );
  Tile mesh_6_6 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177985.4]
    .clock(mesh_6_6_clock),
    .io_in_a_0(mesh_6_6_io_in_a_0),
    .io_in_b_0(mesh_6_6_io_in_b_0),
    .io_in_d_0(mesh_6_6_io_in_d_0),
    .io_in_control_0_propagate(mesh_6_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_6_io_in_control_0_shift),
    .io_out_a_0(mesh_6_6_io_out_a_0),
    .io_out_c_0(mesh_6_6_io_out_c_0),
    .io_out_b_0(mesh_6_6_io_out_b_0),
    .io_out_control_0_propagate(mesh_6_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_6_io_out_control_0_shift),
    .io_in_valid_0(mesh_6_6_io_in_valid_0),
    .io_out_valid_0(mesh_6_6_io_out_valid_0)
  );
  Tile mesh_6_7 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177988.4]
    .clock(mesh_6_7_clock),
    .io_in_a_0(mesh_6_7_io_in_a_0),
    .io_in_b_0(mesh_6_7_io_in_b_0),
    .io_in_d_0(mesh_6_7_io_in_d_0),
    .io_in_control_0_propagate(mesh_6_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_6_7_io_in_control_0_shift),
    .io_out_a_0(mesh_6_7_io_out_a_0),
    .io_out_c_0(mesh_6_7_io_out_c_0),
    .io_out_b_0(mesh_6_7_io_out_b_0),
    .io_out_control_0_propagate(mesh_6_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_6_7_io_out_control_0_shift),
    .io_in_valid_0(mesh_6_7_io_in_valid_0),
    .io_out_valid_0(mesh_6_7_io_out_valid_0)
  );
  Tile mesh_7_0 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177991.4]
    .clock(mesh_7_0_clock),
    .io_in_a_0(mesh_7_0_io_in_a_0),
    .io_in_b_0(mesh_7_0_io_in_b_0),
    .io_in_d_0(mesh_7_0_io_in_d_0),
    .io_in_control_0_propagate(mesh_7_0_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_0_io_in_control_0_shift),
    .io_out_a_0(mesh_7_0_io_out_a_0),
    .io_out_c_0(mesh_7_0_io_out_c_0),
    .io_out_b_0(mesh_7_0_io_out_b_0),
    .io_out_control_0_propagate(mesh_7_0_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_0_io_out_control_0_shift),
    .io_in_valid_0(mesh_7_0_io_in_valid_0),
    .io_out_valid_0(mesh_7_0_io_out_valid_0)
  );
  Tile mesh_7_1 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177994.4]
    .clock(mesh_7_1_clock),
    .io_in_a_0(mesh_7_1_io_in_a_0),
    .io_in_b_0(mesh_7_1_io_in_b_0),
    .io_in_d_0(mesh_7_1_io_in_d_0),
    .io_in_control_0_propagate(mesh_7_1_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_1_io_in_control_0_shift),
    .io_out_a_0(mesh_7_1_io_out_a_0),
    .io_out_c_0(mesh_7_1_io_out_c_0),
    .io_out_b_0(mesh_7_1_io_out_b_0),
    .io_out_control_0_propagate(mesh_7_1_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_1_io_out_control_0_shift),
    .io_in_valid_0(mesh_7_1_io_in_valid_0),
    .io_out_valid_0(mesh_7_1_io_out_valid_0)
  );
  Tile mesh_7_2 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177997.4]
    .clock(mesh_7_2_clock),
    .io_in_a_0(mesh_7_2_io_in_a_0),
    .io_in_b_0(mesh_7_2_io_in_b_0),
    .io_in_d_0(mesh_7_2_io_in_d_0),
    .io_in_control_0_propagate(mesh_7_2_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_2_io_in_control_0_shift),
    .io_out_a_0(mesh_7_2_io_out_a_0),
    .io_out_c_0(mesh_7_2_io_out_c_0),
    .io_out_b_0(mesh_7_2_io_out_b_0),
    .io_out_control_0_propagate(mesh_7_2_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_2_io_out_control_0_shift),
    .io_in_valid_0(mesh_7_2_io_in_valid_0),
    .io_out_valid_0(mesh_7_2_io_out_valid_0)
  );
  Tile mesh_7_3 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178000.4]
    .clock(mesh_7_3_clock),
    .io_in_a_0(mesh_7_3_io_in_a_0),
    .io_in_b_0(mesh_7_3_io_in_b_0),
    .io_in_d_0(mesh_7_3_io_in_d_0),
    .io_in_control_0_propagate(mesh_7_3_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_3_io_in_control_0_shift),
    .io_out_a_0(mesh_7_3_io_out_a_0),
    .io_out_c_0(mesh_7_3_io_out_c_0),
    .io_out_b_0(mesh_7_3_io_out_b_0),
    .io_out_control_0_propagate(mesh_7_3_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_3_io_out_control_0_shift),
    .io_in_valid_0(mesh_7_3_io_in_valid_0),
    .io_out_valid_0(mesh_7_3_io_out_valid_0)
  );
  Tile mesh_7_4 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178003.4]
    .clock(mesh_7_4_clock),
    .io_in_a_0(mesh_7_4_io_in_a_0),
    .io_in_b_0(mesh_7_4_io_in_b_0),
    .io_in_d_0(mesh_7_4_io_in_d_0),
    .io_in_control_0_propagate(mesh_7_4_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_4_io_in_control_0_shift),
    .io_out_a_0(mesh_7_4_io_out_a_0),
    .io_out_c_0(mesh_7_4_io_out_c_0),
    .io_out_b_0(mesh_7_4_io_out_b_0),
    .io_out_control_0_propagate(mesh_7_4_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_4_io_out_control_0_shift),
    .io_in_valid_0(mesh_7_4_io_in_valid_0),
    .io_out_valid_0(mesh_7_4_io_out_valid_0)
  );
  Tile mesh_7_5 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178006.4]
    .clock(mesh_7_5_clock),
    .io_in_a_0(mesh_7_5_io_in_a_0),
    .io_in_b_0(mesh_7_5_io_in_b_0),
    .io_in_d_0(mesh_7_5_io_in_d_0),
    .io_in_control_0_propagate(mesh_7_5_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_5_io_in_control_0_shift),
    .io_out_a_0(mesh_7_5_io_out_a_0),
    .io_out_c_0(mesh_7_5_io_out_c_0),
    .io_out_b_0(mesh_7_5_io_out_b_0),
    .io_out_control_0_propagate(mesh_7_5_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_5_io_out_control_0_shift),
    .io_in_valid_0(mesh_7_5_io_in_valid_0),
    .io_out_valid_0(mesh_7_5_io_out_valid_0)
  );
  Tile mesh_7_6 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178009.4]
    .clock(mesh_7_6_clock),
    .io_in_a_0(mesh_7_6_io_in_a_0),
    .io_in_b_0(mesh_7_6_io_in_b_0),
    .io_in_d_0(mesh_7_6_io_in_d_0),
    .io_in_control_0_propagate(mesh_7_6_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_6_io_in_control_0_shift),
    .io_out_a_0(mesh_7_6_io_out_a_0),
    .io_out_c_0(mesh_7_6_io_out_c_0),
    .io_out_b_0(mesh_7_6_io_out_b_0),
    .io_out_control_0_propagate(mesh_7_6_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_6_io_out_control_0_shift),
    .io_in_valid_0(mesh_7_6_io_in_valid_0),
    .io_out_valid_0(mesh_7_6_io_out_valid_0)
  );
  Tile mesh_7_7 ( // @[Mesh.scala 33:71:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178012.4]
    .clock(mesh_7_7_clock),
    .io_in_a_0(mesh_7_7_io_in_a_0),
    .io_in_b_0(mesh_7_7_io_in_b_0),
    .io_in_d_0(mesh_7_7_io_in_d_0),
    .io_in_control_0_propagate(mesh_7_7_io_in_control_0_propagate),
    .io_in_control_0_shift(mesh_7_7_io_in_control_0_shift),
    .io_out_a_0(mesh_7_7_io_out_a_0),
    .io_out_c_0(mesh_7_7_io_out_c_0),
    .io_out_b_0(mesh_7_7_io_out_b_0),
    .io_out_control_0_propagate(mesh_7_7_io_out_control_0_propagate),
    .io_out_control_0_shift(mesh_7_7_io_out_control_0_shift),
    .io_in_valid_0(mesh_7_7_io_in_valid_0),
    .io_out_valid_0(mesh_7_7_io_out_valid_0)
  );
  
  reg [18:0] _RAND_c00;
reg [64:0] _RAND_b00;

reg [acc_wl-1:0] temp_io_out_c_0_0 ;
reg [acc_wl-1:0] temp_io_out_c_1_0 ;
reg [acc_wl-1:0] temp_io_out_c_2_0 ;
reg [acc_wl-1:0] temp_io_out_c_3_0 ;
reg [acc_wl-1:0] temp_io_out_c_4_0 ;
reg [acc_wl-1:0] temp_io_out_c_5_0 ;
reg [acc_wl-1:0] temp_io_out_c_6_0 ;
reg [acc_wl-1:0] temp_io_out_c_7_0 ;

  
  initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_c00 = {1{`RANDOM}};
  
io_out_c_0_0= _RAND_c00;
io_out_c_1_0= _RAND_c00;
io_out_c_2_0= _RAND_c00;
io_out_c_3_0= _RAND_c00;
io_out_c_4_0= _RAND_c00;
io_out_c_5_0= _RAND_c00;
io_out_c_6_0= _RAND_c00;
io_out_c_7_0= _RAND_c00;
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
_RAND_b00 ={1{`RANDOM}};
temp_io_out_c_0_0=_RAND_b00;
temp_io_out_c_1_0=_RAND_b00;
temp_io_out_c_2_0=_RAND_b00;
temp_io_out_c_3_0=_RAND_b00;
temp_io_out_c_4_0=_RAND_b00;
temp_io_out_c_5_0=_RAND_b00;
temp_io_out_c_6_0=_RAND_b00;
temp_io_out_c_7_0=_RAND_b00;
io_out_valid_0_0=_RAND_b00[0:0];
  
  
  
  
    `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  
always@(posedge clock) begin
temp_io_out_c_0_0 <= {{$signed(mesh_7_0_io_out_c_0[(2*(acc_wl-k)+k-1):acc_wl])+$signed(mesh_7_0_io_out_c_0[acc_wl-1:k])},mesh_7_0_io_out_c_0[k-1:0]};
temp_io_out_c_1_0 <= {{$signed(mesh_7_1_io_out_c_0[(2*(acc_wl-k)+k-1):acc_wl])+$signed(mesh_7_1_io_out_c_0[acc_wl-1:k])},mesh_7_1_io_out_c_0[k-1:0]};
temp_io_out_c_2_0 <= {{$signed(mesh_7_2_io_out_c_0[(2*(acc_wl-k)+k-1):acc_wl])+$signed(mesh_7_2_io_out_c_0[acc_wl-1:k])},mesh_7_2_io_out_c_0[k-1:0]};
temp_io_out_c_3_0 <= {{$signed(mesh_7_3_io_out_c_0[(2*(acc_wl-k)+k-1):acc_wl])+$signed(mesh_7_3_io_out_c_0[acc_wl-1:k])},mesh_7_3_io_out_c_0[k-1:0]};
temp_io_out_c_4_0 <= {{$signed(mesh_7_4_io_out_c_0[(2*(acc_wl-k)+k-1):acc_wl])+$signed(mesh_7_4_io_out_c_0[acc_wl-1:k])},mesh_7_4_io_out_c_0[k-1:0]};
temp_io_out_c_5_0 <= {{$signed(mesh_7_5_io_out_c_0[(2*(acc_wl-k)+k-1):acc_wl])+$signed(mesh_7_5_io_out_c_0[acc_wl-1:k])},mesh_7_5_io_out_c_0[k-1:0]};
temp_io_out_c_6_0 <= {{$signed(mesh_7_6_io_out_c_0[(2*(acc_wl-k)+k-1):acc_wl])+$signed(mesh_7_6_io_out_c_0[acc_wl-1:k])},mesh_7_6_io_out_c_0[k-1:0]};
temp_io_out_c_7_0 <= {{$signed(mesh_7_7_io_out_c_0[(2*(acc_wl-k)+k-1):acc_wl])+$signed(mesh_7_7_io_out_c_0[acc_wl-1:k])},mesh_7_7_io_out_c_0[k-1:0]};
end
wire [18:0] temp_mesh_7_0_io_out_c_0;
wire [18:0] temp_mesh_7_1_io_out_c_0;
wire [18:0] temp_mesh_7_2_io_out_c_0;
wire [18:0] temp_mesh_7_3_io_out_c_0;
wire [18:0] temp_mesh_7_4_io_out_c_0;
wire [18:0] temp_mesh_7_5_io_out_c_0;
wire [18:0] temp_mesh_7_6_io_out_c_0;
wire [18:0] temp_mesh_7_7_io_out_c_0;

rounding round_0(.clock(clock),.c1(temp_io_out_c_0_0),.io_in_control_shift(mesh_7_0_io_out_c_0[(2*(acc_wl-k)+k+5):(2*(acc_wl-k)+k)]),.io_in_control_propagate(mesh_7_0_io_out_c_0[(2*(acc_wl-k)+k+6)]),.io_in_valid(mesh_7_0_io_out_c_0[(2*(acc_wl-k)+k+7)]), ._T_35(temp_mesh_7_0_io_out_c_0));
rounding round_1(.clock(clock),.c1(temp_io_out_c_1_0),.io_in_control_shift(mesh_7_1_io_out_c_0[(2*(acc_wl-k)+k+5):(2*(acc_wl-k)+k)]),.io_in_control_propagate(mesh_7_1_io_out_c_0[(2*(acc_wl-k)+k+6)]),.io_in_valid(mesh_7_1_io_out_c_0[(2*(acc_wl-k)+k+7)]), ._T_35(temp_mesh_7_1_io_out_c_0));
rounding round_2(.clock(clock),.c1(temp_io_out_c_2_0),.io_in_control_shift(mesh_7_2_io_out_c_0[(2*(acc_wl-k)+k+5):(2*(acc_wl-k)+k)]),.io_in_control_propagate(mesh_7_2_io_out_c_0[(2*(acc_wl-k)+k+6)]),.io_in_valid(mesh_7_2_io_out_c_0[(2*(acc_wl-k)+k+7)]), ._T_35(temp_mesh_7_2_io_out_c_0));
rounding round_3(.clock(clock),.c1(temp_io_out_c_3_0),.io_in_control_shift(mesh_7_3_io_out_c_0[(2*(acc_wl-k)+k+5):(2*(acc_wl-k)+k)]),.io_in_control_propagate(mesh_7_3_io_out_c_0[(2*(acc_wl-k)+k+6)]),.io_in_valid(mesh_7_3_io_out_c_0[(2*(acc_wl-k)+k+7)]), ._T_35(temp_mesh_7_3_io_out_c_0));
rounding round_4(.clock(clock),.c1(temp_io_out_c_4_0),.io_in_control_shift(mesh_7_4_io_out_c_0[(2*(acc_wl-k)+k+5):(2*(acc_wl-k)+k)]),.io_in_control_propagate(mesh_7_4_io_out_c_0[(2*(acc_wl-k)+k+6)]),.io_in_valid(mesh_7_4_io_out_c_0[(2*(acc_wl-k)+k+7)]), ._T_35(temp_mesh_7_4_io_out_c_0));
rounding round_5(.clock(clock),.c1(temp_io_out_c_5_0),.io_in_control_shift(mesh_7_5_io_out_c_0[(2*(acc_wl-k)+k+5):(2*(acc_wl-k)+k)]),.io_in_control_propagate(mesh_7_5_io_out_c_0[(2*(acc_wl-k)+k+6)]),.io_in_valid(mesh_7_5_io_out_c_0[(2*(acc_wl-k)+k+7)]), ._T_35(temp_mesh_7_5_io_out_c_0));
rounding round_6(.clock(clock),.c1(temp_io_out_c_6_0),.io_in_control_shift(mesh_7_6_io_out_c_0[(2*(acc_wl-k)+k+5):(2*(acc_wl-k)+k)]),.io_in_control_propagate(mesh_7_6_io_out_c_0[(2*(acc_wl-k)+k+6)]),.io_in_valid(mesh_7_6_io_out_c_0[(2*(acc_wl-k)+k+7)]), ._T_35(temp_mesh_7_6_io_out_c_0));
rounding round_7(.clock(clock),.c1(temp_io_out_c_7_0),.io_in_control_shift(mesh_7_7_io_out_c_0[(2*(acc_wl-k)+k+5):(2*(acc_wl-k)+k)]),.io_in_control_propagate(mesh_7_7_io_out_c_0[(2*(acc_wl-k)+k+6)]),.io_in_valid(mesh_7_7_io_out_c_0[(2*(acc_wl-k)+k+7)]), ._T_35(temp_mesh_7_7_io_out_c_0));

assign io_out_b_0_0 = $signed(temp_mesh_7_0_io_out_c_0);
assign io_out_b_1_0 = $signed(temp_mesh_7_1_io_out_c_0);
assign io_out_b_2_0 = $signed(temp_mesh_7_2_io_out_c_0);
assign io_out_b_3_0 = $signed(temp_mesh_7_3_io_out_c_0);
assign io_out_b_4_0 = $signed(temp_mesh_7_4_io_out_c_0);
assign io_out_b_5_0 = $signed(temp_mesh_7_5_io_out_c_0);
assign io_out_b_6_0 = $signed(temp_mesh_7_6_io_out_c_0);
assign io_out_b_7_0 = $signed(temp_mesh_7_7_io_out_c_0);

always@(posedge clock) begin
io_out_c_0_0 <= mesh_7_0_io_out_b_0;
io_out_c_1_0 <= mesh_7_1_io_out_b_0;
io_out_c_2_0 <= mesh_7_2_io_out_b_0;
io_out_c_3_0 <= mesh_7_3_io_out_b_0;
io_out_c_4_0 <= mesh_7_4_io_out_b_0;
io_out_c_5_0 <= mesh_7_5_io_out_b_0;
io_out_c_6_0 <= mesh_7_6_io_out_b_0;
io_out_c_7_0 <= mesh_7_7_io_out_b_0;
io_out_valid_0_0 <= mesh_7_0_io_out_valid_0;
end
  
  
  
  //assign io_out_c_0_0 = mesh_7_0_io_out_b_0; // @[Mesh.scala 85:7:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180143.4]
  //assign io_out_c_1_0 = mesh_7_1_io_out_b_0; // @[Mesh.scala 85:7:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180146.4]
  //assign io_out_c_2_0 = mesh_7_2_io_out_b_0; // @[Mesh.scala 85:7:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180149.4]
  //assign io_out_c_3_0 = mesh_7_3_io_out_b_0; // @[Mesh.scala 85:7:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180152.4]
  //assign io_out_c_4_0 = mesh_7_4_io_out_b_0; // @[Mesh.scala 85:7:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180155.4]
  //assign io_out_c_5_0 = mesh_7_5_io_out_b_0; // @[Mesh.scala 85:7:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180158.4]
  //assign io_out_c_6_0 = mesh_7_6_io_out_b_0; // @[Mesh.scala 85:7:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180161.4]
  //assign io_out_c_7_0 = mesh_7_7_io_out_b_0; // @[Mesh.scala 85:7:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180164.4]
  //assign io_out_b_0_0 = mesh_7_0_io_out_c_0; // @[Mesh.scala 86:7:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180144.4]
  //assign io_out_b_1_0 = mesh_7_1_io_out_c_0; // @[Mesh.scala 86:7:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180147.4]
  //assign io_out_b_2_0 = mesh_7_2_io_out_c_0; // @[Mesh.scala 86:7:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180150.4]
  //assign io_out_b_3_0 = mesh_7_3_io_out_c_0; // @[Mesh.scala 86:7:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180153.4]
  //assign io_out_b_4_0 = mesh_7_4_io_out_c_0; // @[Mesh.scala 86:7:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180156.4]
  //assign io_out_b_5_0 = mesh_7_5_io_out_c_0; // @[Mesh.scala 86:7:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180159.4]
  //assign io_out_b_6_0 = mesh_7_6_io_out_c_0; // @[Mesh.scala 86:7:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180162.4]
  //assign io_out_b_7_0 = mesh_7_7_io_out_c_0; // @[Mesh.scala 86:7:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180165.4]
  //assign io_out_valid_0_0 = mesh_7_0_io_out_valid_0; // @[Mesh.scala 87:7:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180145.4]
  
  assign mesh_0_0_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177824.4]
  assign mesh_0_0_io_in_a_0 = _T_1_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178019.4]
  assign mesh_0_0_io_in_b_0 = {{11{_T_74_0[7]}},_T_74_0}; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178231.4]
  assign mesh_0_0_io_in_d_0 = {{11{_T_154_0[7]}},_T_154_0}; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178583.4]
  assign mesh_0_0_io_in_control_0_propagate = _T_236; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178947.4]
  assign mesh_0_0_io_in_control_0_shift = _T_234; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178937.4]
  assign mesh_0_0_io_in_valid_0 = _T_441_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179939.4]
  assign mesh_0_1_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177827.4]
  assign mesh_0_1_io_in_a_0 = _T_2_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178022.4]
  assign mesh_0_1_io_in_b_0 = {{11{_T_84_0[7]}},_T_84_0}; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178275.4]
  assign mesh_0_1_io_in_d_0 = {{11{_T_164_0[7]}},_T_164_0}; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178627.4]
  assign mesh_0_1_io_in_control_0_propagate = _T_262; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179073.4]
  assign mesh_0_1_io_in_control_0_shift = _T_260; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179063.4]
  assign mesh_0_1_io_in_valid_0 = _T_450_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179965.4]
  assign mesh_0_2_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177830.4]
  assign mesh_0_2_io_in_a_0 = _T_3_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178025.4]
  assign mesh_0_2_io_in_b_0 = {{11{_T_94_0[7]}},_T_94_0}; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178319.4]
  assign mesh_0_2_io_in_d_0 = {{11{_T_174_0[7]}},_T_174_0}; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178671.4]
  assign mesh_0_2_io_in_control_0_propagate = _T_288; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179199.4]
  assign mesh_0_2_io_in_control_0_shift = _T_286; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179189.4]
  assign mesh_0_2_io_in_valid_0 = _T_459_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179991.4]
  assign mesh_0_3_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177833.4]
  assign mesh_0_3_io_in_a_0 = _T_4_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178028.4]
  assign mesh_0_3_io_in_b_0 = {{11{_T_104_0[7]}},_T_104_0}; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178363.4]
  assign mesh_0_3_io_in_d_0 = {{11{_T_184_0[7]}},_T_184_0}; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178715.4]
  assign mesh_0_3_io_in_control_0_propagate = _T_314; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179325.4]
  assign mesh_0_3_io_in_control_0_shift = _T_312; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179315.4]
  assign mesh_0_3_io_in_valid_0 = _T_468_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180017.4]
  assign mesh_0_4_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177836.4]
  assign mesh_0_4_io_in_a_0 = _T_5_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178031.4]
  assign mesh_0_4_io_in_b_0 = {{11{_T_114_0[7]}},_T_114_0}; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178407.4]
  assign mesh_0_4_io_in_d_0 = {{11{_T_194_0[7]}},_T_194_0}; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178759.4]
  assign mesh_0_4_io_in_control_0_propagate = _T_340; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179451.4]
  assign mesh_0_4_io_in_control_0_shift = _T_338; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179441.4]
  assign mesh_0_4_io_in_valid_0 = _T_477_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180043.4]
  assign mesh_0_5_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177839.4]
  assign mesh_0_5_io_in_a_0 = _T_6_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178034.4]
  assign mesh_0_5_io_in_b_0 = {{11{_T_124_0[7]}},_T_124_0}; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178451.4]
  assign mesh_0_5_io_in_d_0 = {{11{_T_204_0[7]}},_T_204_0}; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178803.4]
  assign mesh_0_5_io_in_control_0_propagate = _T_366; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179577.4]
  assign mesh_0_5_io_in_control_0_shift = _T_364; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179567.4]
  assign mesh_0_5_io_in_valid_0 = _T_486_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180069.4]
  assign mesh_0_6_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177842.4]
  assign mesh_0_6_io_in_a_0 = _T_7_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178037.4]
  assign mesh_0_6_io_in_b_0 = {{11{_T_134_0[7]}},_T_134_0}; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178495.4]
  assign mesh_0_6_io_in_d_0 = {{11{_T_214_0[7]}},_T_214_0}; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178847.4]
  assign mesh_0_6_io_in_control_0_propagate = _T_392; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179703.4]
  assign mesh_0_6_io_in_control_0_shift = _T_390; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179693.4]
  assign mesh_0_6_io_in_valid_0 = _T_495_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180095.4]
  assign mesh_0_7_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177845.4]
  assign mesh_0_7_io_in_a_0 = _T_8_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178040.4]
  assign mesh_0_7_io_in_b_0 = {{11{_T_144_0[7]}},_T_144_0}; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178539.4]
  assign mesh_0_7_io_in_d_0 = {{11{_T_224_0[7]}},_T_224_0}; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178891.4]
  assign mesh_0_7_io_in_control_0_propagate = _T_418; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179829.4]
  assign mesh_0_7_io_in_control_0_shift = _T_416; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179819.4]
  assign mesh_0_7_io_in_valid_0 = _T_504_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180121.4]
  assign mesh_1_0_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177848.4]
  assign mesh_1_0_io_in_a_0 = _T_10_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178045.4]
  assign mesh_1_0_io_in_b_0 = _T_75_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178236.4]
  assign mesh_1_0_io_in_d_0 = _T_155_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178588.4]
  assign mesh_1_0_io_in_control_0_propagate = _T_239; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178962.4]
  assign mesh_1_0_io_in_control_0_shift = _T_237; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178952.4]
  assign mesh_1_0_io_in_valid_0 = _T_442_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179942.4]
  assign mesh_1_1_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177851.4]
  assign mesh_1_1_io_in_a_0 = _T_11_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178048.4]
  assign mesh_1_1_io_in_b_0 = _T_85_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178280.4]
  assign mesh_1_1_io_in_d_0 = _T_165_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178632.4]
  assign mesh_1_1_io_in_control_0_propagate = _T_265; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179088.4]
  assign mesh_1_1_io_in_control_0_shift = _T_263; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179078.4]
  assign mesh_1_1_io_in_valid_0 = _T_451_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179968.4]
  assign mesh_1_2_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177854.4]
  assign mesh_1_2_io_in_a_0 = _T_12_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178051.4]
  assign mesh_1_2_io_in_b_0 = _T_95_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178324.4]
  assign mesh_1_2_io_in_d_0 = _T_175_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178676.4]
  assign mesh_1_2_io_in_control_0_propagate = _T_291; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179214.4]
  assign mesh_1_2_io_in_control_0_shift = _T_289; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179204.4]
  assign mesh_1_2_io_in_valid_0 = _T_460_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179994.4]
  assign mesh_1_3_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177857.4]
  assign mesh_1_3_io_in_a_0 = _T_13_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178054.4]
  assign mesh_1_3_io_in_b_0 = _T_105_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178368.4]
  assign mesh_1_3_io_in_d_0 = _T_185_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178720.4]
  assign mesh_1_3_io_in_control_0_propagate = _T_317; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179340.4]
  assign mesh_1_3_io_in_control_0_shift = _T_315; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179330.4]
  assign mesh_1_3_io_in_valid_0 = _T_469_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180020.4]
  assign mesh_1_4_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177860.4]
  assign mesh_1_4_io_in_a_0 = _T_14_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178057.4]
  assign mesh_1_4_io_in_b_0 = _T_115_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178412.4]
  assign mesh_1_4_io_in_d_0 = _T_195_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178764.4]
  assign mesh_1_4_io_in_control_0_propagate = _T_343; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179466.4]
  assign mesh_1_4_io_in_control_0_shift = _T_341; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179456.4]
  assign mesh_1_4_io_in_valid_0 = _T_478_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180046.4]
  assign mesh_1_5_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177863.4]
  assign mesh_1_5_io_in_a_0 = _T_15_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178060.4]
  assign mesh_1_5_io_in_b_0 = _T_125_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178456.4]
  assign mesh_1_5_io_in_d_0 = _T_205_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178808.4]
  assign mesh_1_5_io_in_control_0_propagate = _T_369; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179592.4]
  assign mesh_1_5_io_in_control_0_shift = _T_367; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179582.4]
  assign mesh_1_5_io_in_valid_0 = _T_487_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180072.4]
  assign mesh_1_6_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177866.4]
  assign mesh_1_6_io_in_a_0 = _T_16_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178063.4]
  assign mesh_1_6_io_in_b_0 = _T_135_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178500.4]
  assign mesh_1_6_io_in_d_0 = _T_215_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178852.4]
  assign mesh_1_6_io_in_control_0_propagate = _T_395; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179718.4]
  assign mesh_1_6_io_in_control_0_shift = _T_393; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179708.4]
  assign mesh_1_6_io_in_valid_0 = _T_496_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180098.4]
  assign mesh_1_7_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177869.4]
  assign mesh_1_7_io_in_a_0 = _T_17_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178066.4]
  assign mesh_1_7_io_in_b_0 = _T_145_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178544.4]
  assign mesh_1_7_io_in_d_0 = _T_225_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178896.4]
  assign mesh_1_7_io_in_control_0_propagate = _T_421; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179844.4]
  assign mesh_1_7_io_in_control_0_shift = _T_419; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179834.4]
  assign mesh_1_7_io_in_valid_0 = _T_505_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180124.4]
  assign mesh_2_0_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177872.4]
  assign mesh_2_0_io_in_a_0 = _T_19_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178071.4]
  assign mesh_2_0_io_in_b_0 = _T_76_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178241.4]
  assign mesh_2_0_io_in_d_0 = _T_156_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178593.4]
  assign mesh_2_0_io_in_control_0_propagate = _T_242; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178977.4]
  assign mesh_2_0_io_in_control_0_shift = _T_240; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178967.4]
  assign mesh_2_0_io_in_valid_0 = _T_443_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179945.4]
  assign mesh_2_1_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177875.4]
  assign mesh_2_1_io_in_a_0 = _T_20_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178074.4]
  assign mesh_2_1_io_in_b_0 = _T_86_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178285.4]
  assign mesh_2_1_io_in_d_0 = _T_166_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178637.4]
  assign mesh_2_1_io_in_control_0_propagate = _T_268; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179103.4]
  assign mesh_2_1_io_in_control_0_shift = _T_266; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179093.4]
  assign mesh_2_1_io_in_valid_0 = _T_452_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179971.4]
  assign mesh_2_2_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177878.4]
  assign mesh_2_2_io_in_a_0 = _T_21_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178077.4]
  assign mesh_2_2_io_in_b_0 = _T_96_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178329.4]
  assign mesh_2_2_io_in_d_0 = _T_176_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178681.4]
  assign mesh_2_2_io_in_control_0_propagate = _T_294; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179229.4]
  assign mesh_2_2_io_in_control_0_shift = _T_292; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179219.4]
  assign mesh_2_2_io_in_valid_0 = _T_461_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179997.4]
  assign mesh_2_3_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177881.4]
  assign mesh_2_3_io_in_a_0 = _T_22_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178080.4]
  assign mesh_2_3_io_in_b_0 = _T_106_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178373.4]
  assign mesh_2_3_io_in_d_0 = _T_186_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178725.4]
  assign mesh_2_3_io_in_control_0_propagate = _T_320; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179355.4]
  assign mesh_2_3_io_in_control_0_shift = _T_318; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179345.4]
  assign mesh_2_3_io_in_valid_0 = _T_470_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180023.4]
  assign mesh_2_4_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177884.4]
  assign mesh_2_4_io_in_a_0 = _T_23_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178083.4]
  assign mesh_2_4_io_in_b_0 = _T_116_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178417.4]
  assign mesh_2_4_io_in_d_0 = _T_196_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178769.4]
  assign mesh_2_4_io_in_control_0_propagate = _T_346; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179481.4]
  assign mesh_2_4_io_in_control_0_shift = _T_344; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179471.4]
  assign mesh_2_4_io_in_valid_0 = _T_479_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180049.4]
  assign mesh_2_5_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177887.4]
  assign mesh_2_5_io_in_a_0 = _T_24_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178086.4]
  assign mesh_2_5_io_in_b_0 = _T_126_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178461.4]
  assign mesh_2_5_io_in_d_0 = _T_206_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178813.4]
  assign mesh_2_5_io_in_control_0_propagate = _T_372; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179607.4]
  assign mesh_2_5_io_in_control_0_shift = _T_370; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179597.4]
  assign mesh_2_5_io_in_valid_0 = _T_488_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180075.4]
  assign mesh_2_6_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177890.4]
  assign mesh_2_6_io_in_a_0 = _T_25_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178089.4]
  assign mesh_2_6_io_in_b_0 = _T_136_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178505.4]
  assign mesh_2_6_io_in_d_0 = _T_216_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178857.4]
  assign mesh_2_6_io_in_control_0_propagate = _T_398; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179733.4]
  assign mesh_2_6_io_in_control_0_shift = _T_396; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179723.4]
  assign mesh_2_6_io_in_valid_0 = _T_497_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180101.4]
  assign mesh_2_7_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177893.4]
  assign mesh_2_7_io_in_a_0 = _T_26_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178092.4]
  assign mesh_2_7_io_in_b_0 = _T_146_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178549.4]
  assign mesh_2_7_io_in_d_0 = _T_226_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178901.4]
  assign mesh_2_7_io_in_control_0_propagate = _T_424; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179859.4]
  assign mesh_2_7_io_in_control_0_shift = _T_422; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179849.4]
  assign mesh_2_7_io_in_valid_0 = _T_506_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180127.4]
  assign mesh_3_0_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177896.4]
  assign mesh_3_0_io_in_a_0 = _T_28_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178097.4]
  assign mesh_3_0_io_in_b_0 = _T_77_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178246.4]
  assign mesh_3_0_io_in_d_0 = _T_157_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178598.4]
  assign mesh_3_0_io_in_control_0_propagate = _T_245; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178992.4]
  assign mesh_3_0_io_in_control_0_shift = _T_243; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178982.4]
  assign mesh_3_0_io_in_valid_0 = _T_444_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179948.4]
  assign mesh_3_1_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177899.4]
  assign mesh_3_1_io_in_a_0 = _T_29_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178100.4]
  assign mesh_3_1_io_in_b_0 = _T_87_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178290.4]
  assign mesh_3_1_io_in_d_0 = _T_167_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178642.4]
  assign mesh_3_1_io_in_control_0_propagate = _T_271; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179118.4]
  assign mesh_3_1_io_in_control_0_shift = _T_269; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179108.4]
  assign mesh_3_1_io_in_valid_0 = _T_453_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179974.4]
  assign mesh_3_2_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177902.4]
  assign mesh_3_2_io_in_a_0 = _T_30_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178103.4]
  assign mesh_3_2_io_in_b_0 = _T_97_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178334.4]
  assign mesh_3_2_io_in_d_0 = _T_177_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178686.4]
  assign mesh_3_2_io_in_control_0_propagate = _T_297; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179244.4]
  assign mesh_3_2_io_in_control_0_shift = _T_295; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179234.4]
  assign mesh_3_2_io_in_valid_0 = _T_462_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180000.4]
  assign mesh_3_3_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177905.4]
  assign mesh_3_3_io_in_a_0 = _T_31_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178106.4]
  assign mesh_3_3_io_in_b_0 = _T_107_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178378.4]
  assign mesh_3_3_io_in_d_0 = _T_187_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178730.4]
  assign mesh_3_3_io_in_control_0_propagate = _T_323; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179370.4]
  assign mesh_3_3_io_in_control_0_shift = _T_321; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179360.4]
  assign mesh_3_3_io_in_valid_0 = _T_471_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180026.4]
  assign mesh_3_4_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177908.4]
  assign mesh_3_4_io_in_a_0 = _T_32_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178109.4]
  assign mesh_3_4_io_in_b_0 = _T_117_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178422.4]
  assign mesh_3_4_io_in_d_0 = _T_197_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178774.4]
  assign mesh_3_4_io_in_control_0_propagate = _T_349; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179496.4]
  assign mesh_3_4_io_in_control_0_shift = _T_347; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179486.4]
  assign mesh_3_4_io_in_valid_0 = _T_480_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180052.4]
  assign mesh_3_5_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177911.4]
  assign mesh_3_5_io_in_a_0 = _T_33_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178112.4]
  assign mesh_3_5_io_in_b_0 = _T_127_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178466.4]
  assign mesh_3_5_io_in_d_0 = _T_207_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178818.4]
  assign mesh_3_5_io_in_control_0_propagate = _T_375; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179622.4]
  assign mesh_3_5_io_in_control_0_shift = _T_373; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179612.4]
  assign mesh_3_5_io_in_valid_0 = _T_489_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180078.4]
  assign mesh_3_6_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177914.4]
  assign mesh_3_6_io_in_a_0 = _T_34_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178115.4]
  assign mesh_3_6_io_in_b_0 = _T_137_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178510.4]
  assign mesh_3_6_io_in_d_0 = _T_217_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178862.4]
  assign mesh_3_6_io_in_control_0_propagate = _T_401; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179748.4]
  assign mesh_3_6_io_in_control_0_shift = _T_399; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179738.4]
  assign mesh_3_6_io_in_valid_0 = _T_498_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180104.4]
  assign mesh_3_7_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177917.4]
  assign mesh_3_7_io_in_a_0 = _T_35_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178118.4]
  assign mesh_3_7_io_in_b_0 = _T_147_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178554.4]
  assign mesh_3_7_io_in_d_0 = _T_227_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178906.4]
  assign mesh_3_7_io_in_control_0_propagate = _T_427; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179874.4]
  assign mesh_3_7_io_in_control_0_shift = _T_425; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179864.4]
  assign mesh_3_7_io_in_valid_0 = _T_507_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180130.4]
  assign mesh_4_0_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177920.4]
  assign mesh_4_0_io_in_a_0 = _T_37_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178123.4]
  assign mesh_4_0_io_in_b_0 = _T_78_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178251.4]
  assign mesh_4_0_io_in_d_0 = _T_158_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178603.4]
  assign mesh_4_0_io_in_control_0_propagate = _T_248; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179007.4]
  assign mesh_4_0_io_in_control_0_shift = _T_246; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178997.4]
  assign mesh_4_0_io_in_valid_0 = _T_445_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179951.4]
  assign mesh_4_1_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177923.4]
  assign mesh_4_1_io_in_a_0 = _T_38_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178126.4]
  assign mesh_4_1_io_in_b_0 = _T_88_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178295.4]
  assign mesh_4_1_io_in_d_0 = _T_168_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178647.4]
  assign mesh_4_1_io_in_control_0_propagate = _T_274; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179133.4]
  assign mesh_4_1_io_in_control_0_shift = _T_272; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179123.4]
  assign mesh_4_1_io_in_valid_0 = _T_454_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179977.4]
  assign mesh_4_2_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177926.4]
  assign mesh_4_2_io_in_a_0 = _T_39_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178129.4]
  assign mesh_4_2_io_in_b_0 = _T_98_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178339.4]
  assign mesh_4_2_io_in_d_0 = _T_178_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178691.4]
  assign mesh_4_2_io_in_control_0_propagate = _T_300; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179259.4]
  assign mesh_4_2_io_in_control_0_shift = _T_298; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179249.4]
  assign mesh_4_2_io_in_valid_0 = _T_463_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180003.4]
  assign mesh_4_3_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177929.4]
  assign mesh_4_3_io_in_a_0 = _T_40_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178132.4]
  assign mesh_4_3_io_in_b_0 = _T_108_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178383.4]
  assign mesh_4_3_io_in_d_0 = _T_188_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178735.4]
  assign mesh_4_3_io_in_control_0_propagate = _T_326; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179385.4]
  assign mesh_4_3_io_in_control_0_shift = _T_324; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179375.4]
  assign mesh_4_3_io_in_valid_0 = _T_472_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180029.4]
  assign mesh_4_4_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177932.4]
  assign mesh_4_4_io_in_a_0 = _T_41_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178135.4]
  assign mesh_4_4_io_in_b_0 = _T_118_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178427.4]
  assign mesh_4_4_io_in_d_0 = _T_198_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178779.4]
  assign mesh_4_4_io_in_control_0_propagate = _T_352; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179511.4]
  assign mesh_4_4_io_in_control_0_shift = _T_350; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179501.4]
  assign mesh_4_4_io_in_valid_0 = _T_481_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180055.4]
  assign mesh_4_5_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177935.4]
  assign mesh_4_5_io_in_a_0 = _T_42_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178138.4]
  assign mesh_4_5_io_in_b_0 = _T_128_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178471.4]
  assign mesh_4_5_io_in_d_0 = _T_208_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178823.4]
  assign mesh_4_5_io_in_control_0_propagate = _T_378; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179637.4]
  assign mesh_4_5_io_in_control_0_shift = _T_376; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179627.4]
  assign mesh_4_5_io_in_valid_0 = _T_490_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180081.4]
  assign mesh_4_6_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177938.4]
  assign mesh_4_6_io_in_a_0 = _T_43_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178141.4]
  assign mesh_4_6_io_in_b_0 = _T_138_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178515.4]
  assign mesh_4_6_io_in_d_0 = _T_218_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178867.4]
  assign mesh_4_6_io_in_control_0_propagate = _T_404; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179763.4]
  assign mesh_4_6_io_in_control_0_shift = _T_402; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179753.4]
  assign mesh_4_6_io_in_valid_0 = _T_499_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180107.4]
  assign mesh_4_7_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177941.4]
  assign mesh_4_7_io_in_a_0 = _T_44_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178144.4]
  assign mesh_4_7_io_in_b_0 = _T_148_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178559.4]
  assign mesh_4_7_io_in_d_0 = _T_228_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178911.4]
  assign mesh_4_7_io_in_control_0_propagate = _T_430; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179889.4]
  assign mesh_4_7_io_in_control_0_shift = _T_428; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179879.4]
  assign mesh_4_7_io_in_valid_0 = _T_508_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180133.4]
  assign mesh_5_0_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177944.4]
  assign mesh_5_0_io_in_a_0 = _T_46_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178149.4]
  assign mesh_5_0_io_in_b_0 = _T_79_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178256.4]
  assign mesh_5_0_io_in_d_0 = _T_159_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178608.4]
  assign mesh_5_0_io_in_control_0_propagate = _T_251; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179022.4]
  assign mesh_5_0_io_in_control_0_shift = _T_249; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179012.4]
  assign mesh_5_0_io_in_valid_0 = _T_446_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179954.4]
  assign mesh_5_1_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177947.4]
  assign mesh_5_1_io_in_a_0 = _T_47_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178152.4]
  assign mesh_5_1_io_in_b_0 = _T_89_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178300.4]
  assign mesh_5_1_io_in_d_0 = _T_169_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178652.4]
  assign mesh_5_1_io_in_control_0_propagate = _T_277; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179148.4]
  assign mesh_5_1_io_in_control_0_shift = _T_275; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179138.4]
  assign mesh_5_1_io_in_valid_0 = _T_455_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179980.4]
  assign mesh_5_2_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177950.4]
  assign mesh_5_2_io_in_a_0 = _T_48_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178155.4]
  assign mesh_5_2_io_in_b_0 = _T_99_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178344.4]
  assign mesh_5_2_io_in_d_0 = _T_179_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178696.4]
  assign mesh_5_2_io_in_control_0_propagate = _T_303; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179274.4]
  assign mesh_5_2_io_in_control_0_shift = _T_301; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179264.4]
  assign mesh_5_2_io_in_valid_0 = _T_464_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180006.4]
  assign mesh_5_3_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177953.4]
  assign mesh_5_3_io_in_a_0 = _T_49_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178158.4]
  assign mesh_5_3_io_in_b_0 = _T_109_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178388.4]
  assign mesh_5_3_io_in_d_0 = _T_189_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178740.4]
  assign mesh_5_3_io_in_control_0_propagate = _T_329; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179400.4]
  assign mesh_5_3_io_in_control_0_shift = _T_327; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179390.4]
  assign mesh_5_3_io_in_valid_0 = _T_473_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180032.4]
  assign mesh_5_4_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177956.4]
  assign mesh_5_4_io_in_a_0 = _T_50_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178161.4]
  assign mesh_5_4_io_in_b_0 = _T_119_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178432.4]
  assign mesh_5_4_io_in_d_0 = _T_199_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178784.4]
  assign mesh_5_4_io_in_control_0_propagate = _T_355; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179526.4]
  assign mesh_5_4_io_in_control_0_shift = _T_353; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179516.4]
  assign mesh_5_4_io_in_valid_0 = _T_482_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180058.4]
  assign mesh_5_5_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177959.4]
  assign mesh_5_5_io_in_a_0 = _T_51_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178164.4]
  assign mesh_5_5_io_in_b_0 = _T_129_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178476.4]
  assign mesh_5_5_io_in_d_0 = _T_209_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178828.4]
  assign mesh_5_5_io_in_control_0_propagate = _T_381; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179652.4]
  assign mesh_5_5_io_in_control_0_shift = _T_379; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179642.4]
  assign mesh_5_5_io_in_valid_0 = _T_491_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180084.4]
  assign mesh_5_6_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177962.4]
  assign mesh_5_6_io_in_a_0 = _T_52_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178167.4]
  assign mesh_5_6_io_in_b_0 = _T_139_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178520.4]
  assign mesh_5_6_io_in_d_0 = _T_219_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178872.4]
  assign mesh_5_6_io_in_control_0_propagate = _T_407; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179778.4]
  assign mesh_5_6_io_in_control_0_shift = _T_405; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179768.4]
  assign mesh_5_6_io_in_valid_0 = _T_500_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180110.4]
  assign mesh_5_7_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177965.4]
  assign mesh_5_7_io_in_a_0 = _T_53_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178170.4]
  assign mesh_5_7_io_in_b_0 = _T_149_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178564.4]
  assign mesh_5_7_io_in_d_0 = _T_229_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178916.4]
  assign mesh_5_7_io_in_control_0_propagate = _T_433; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179904.4]
  assign mesh_5_7_io_in_control_0_shift = _T_431; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179894.4]
  assign mesh_5_7_io_in_valid_0 = _T_509_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180136.4]
  assign mesh_6_0_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177968.4]
  assign mesh_6_0_io_in_a_0 = _T_55_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178175.4]
  assign mesh_6_0_io_in_b_0 = _T_80_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178261.4]
  assign mesh_6_0_io_in_d_0 = _T_160_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178613.4]
  assign mesh_6_0_io_in_control_0_propagate = _T_254; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179037.4]
  assign mesh_6_0_io_in_control_0_shift = _T_252; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179027.4]
  assign mesh_6_0_io_in_valid_0 = _T_447_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179957.4]
  assign mesh_6_1_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177971.4]
  assign mesh_6_1_io_in_a_0 = _T_56_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178178.4]
  assign mesh_6_1_io_in_b_0 = _T_90_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178305.4]
  assign mesh_6_1_io_in_d_0 = _T_170_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178657.4]
  assign mesh_6_1_io_in_control_0_propagate = _T_280; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179163.4]
  assign mesh_6_1_io_in_control_0_shift = _T_278; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179153.4]
  assign mesh_6_1_io_in_valid_0 = _T_456_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179983.4]
  assign mesh_6_2_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177974.4]
  assign mesh_6_2_io_in_a_0 = _T_57_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178181.4]
  assign mesh_6_2_io_in_b_0 = _T_100_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178349.4]
  assign mesh_6_2_io_in_d_0 = _T_180_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178701.4]
  assign mesh_6_2_io_in_control_0_propagate = _T_306; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179289.4]
  assign mesh_6_2_io_in_control_0_shift = _T_304; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179279.4]
  assign mesh_6_2_io_in_valid_0 = _T_465_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180009.4]
  assign mesh_6_3_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177977.4]
  assign mesh_6_3_io_in_a_0 = _T_58_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178184.4]
  assign mesh_6_3_io_in_b_0 = _T_110_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178393.4]
  assign mesh_6_3_io_in_d_0 = _T_190_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178745.4]
  assign mesh_6_3_io_in_control_0_propagate = _T_332; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179415.4]
  assign mesh_6_3_io_in_control_0_shift = _T_330; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179405.4]
  assign mesh_6_3_io_in_valid_0 = _T_474_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180035.4]
  assign mesh_6_4_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177980.4]
  assign mesh_6_4_io_in_a_0 = _T_59_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178187.4]
  assign mesh_6_4_io_in_b_0 = _T_120_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178437.4]
  assign mesh_6_4_io_in_d_0 = _T_200_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178789.4]
  assign mesh_6_4_io_in_control_0_propagate = _T_358; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179541.4]
  assign mesh_6_4_io_in_control_0_shift = _T_356; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179531.4]
  assign mesh_6_4_io_in_valid_0 = _T_483_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180061.4]
  assign mesh_6_5_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177983.4]
  assign mesh_6_5_io_in_a_0 = _T_60_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178190.4]
  assign mesh_6_5_io_in_b_0 = _T_130_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178481.4]
  assign mesh_6_5_io_in_d_0 = _T_210_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178833.4]
  assign mesh_6_5_io_in_control_0_propagate = _T_384; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179667.4]
  assign mesh_6_5_io_in_control_0_shift = _T_382; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179657.4]
  assign mesh_6_5_io_in_valid_0 = _T_492_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180087.4]
  assign mesh_6_6_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177986.4]
  assign mesh_6_6_io_in_a_0 = _T_61_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178193.4]
  assign mesh_6_6_io_in_b_0 = _T_140_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178525.4]
  assign mesh_6_6_io_in_d_0 = _T_220_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178877.4]
  assign mesh_6_6_io_in_control_0_propagate = _T_410; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179793.4]
  assign mesh_6_6_io_in_control_0_shift = _T_408; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179783.4]
  assign mesh_6_6_io_in_valid_0 = _T_501_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180113.4]
  assign mesh_6_7_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177989.4]
  assign mesh_6_7_io_in_a_0 = _T_62_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178196.4]
  assign mesh_6_7_io_in_b_0 = _T_150_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178569.4]
  assign mesh_6_7_io_in_d_0 = _T_230_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178921.4]
  assign mesh_6_7_io_in_control_0_propagate = _T_436; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179919.4]
  assign mesh_6_7_io_in_control_0_shift = _T_434; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179909.4]
  assign mesh_6_7_io_in_valid_0 = _T_510_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180139.4]
  assign mesh_7_0_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177992.4]
  assign mesh_7_0_io_in_a_0 = _T_64_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178201.4]
  assign mesh_7_0_io_in_b_0 = _T_81_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178266.4]
  assign mesh_7_0_io_in_d_0 = _T_161_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178618.4]
  assign mesh_7_0_io_in_control_0_propagate = _T_257; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179052.4]
  assign mesh_7_0_io_in_control_0_shift = _T_255; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179042.4]
  assign mesh_7_0_io_in_valid_0 = _T_448_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179960.4]
  assign mesh_7_1_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177995.4]
  assign mesh_7_1_io_in_a_0 = _T_65_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178204.4]
  assign mesh_7_1_io_in_b_0 = _T_91_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178310.4]
  assign mesh_7_1_io_in_d_0 = _T_171_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178662.4]
  assign mesh_7_1_io_in_control_0_propagate = _T_283; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179178.4]
  assign mesh_7_1_io_in_control_0_shift = _T_281; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179168.4]
  assign mesh_7_1_io_in_valid_0 = _T_457_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179986.4]
  assign mesh_7_2_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@177998.4]
  assign mesh_7_2_io_in_a_0 = _T_66_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178207.4]
  assign mesh_7_2_io_in_b_0 = _T_101_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178354.4]
  assign mesh_7_2_io_in_d_0 = _T_181_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178706.4]
  assign mesh_7_2_io_in_control_0_propagate = _T_309; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179304.4]
  assign mesh_7_2_io_in_control_0_shift = _T_307; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179294.4]
  assign mesh_7_2_io_in_valid_0 = _T_466_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180012.4]
  assign mesh_7_3_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178001.4]
  assign mesh_7_3_io_in_a_0 = _T_67_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178210.4]
  assign mesh_7_3_io_in_b_0 = _T_111_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178398.4]
  assign mesh_7_3_io_in_d_0 = _T_191_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178750.4]
  assign mesh_7_3_io_in_control_0_propagate = _T_335; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179430.4]
  assign mesh_7_3_io_in_control_0_shift = _T_333; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179420.4]
  assign mesh_7_3_io_in_valid_0 = _T_475_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180038.4]
  assign mesh_7_4_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178004.4]
  assign mesh_7_4_io_in_a_0 = _T_68_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178213.4]
  assign mesh_7_4_io_in_b_0 = _T_121_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178442.4]
  assign mesh_7_4_io_in_d_0 = _T_201_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178794.4]
  assign mesh_7_4_io_in_control_0_propagate = _T_361; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179556.4]
  assign mesh_7_4_io_in_control_0_shift = _T_359; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179546.4]
  assign mesh_7_4_io_in_valid_0 = _T_484_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180064.4]
  assign mesh_7_5_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178007.4]
  assign mesh_7_5_io_in_a_0 = _T_69_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178216.4]
  assign mesh_7_5_io_in_b_0 = _T_131_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178486.4]
  assign mesh_7_5_io_in_d_0 = _T_211_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178838.4]
  assign mesh_7_5_io_in_control_0_propagate = _T_387; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179682.4]
  assign mesh_7_5_io_in_control_0_shift = _T_385; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179672.4]
  assign mesh_7_5_io_in_valid_0 = _T_493_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180090.4]
  assign mesh_7_6_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178010.4]
  assign mesh_7_6_io_in_a_0 = _T_70_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178219.4]
  assign mesh_7_6_io_in_b_0 = _T_141_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178530.4]
  assign mesh_7_6_io_in_d_0 = _T_221_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178882.4]
  assign mesh_7_6_io_in_control_0_propagate = _T_413; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179808.4]
  assign mesh_7_6_io_in_control_0_shift = _T_411; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179798.4]
  assign mesh_7_6_io_in_valid_0 = _T_502_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180116.4]
  assign mesh_7_7_clock = clock; // @[:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178013.4]
  assign mesh_7_7_io_in_a_0 = _T_71_0; // @[Mesh.scala 42:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178222.4]
  assign mesh_7_7_io_in_b_0 = _T_151_0; // @[Mesh.scala 50:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178574.4]
  assign mesh_7_7_io_in_d_0 = _T_231_0; // @[Mesh.scala 58:22:example.TestHarness.GemminiSocTest1RocketConfig864.fir@178926.4]
  assign mesh_7_7_io_in_control_0_propagate = _T_439; // @[Mesh.scala 69:31:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179934.4]
  assign mesh_7_7_io_in_control_0_shift = _T_437; // @[Mesh.scala 67:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@179924.4]
  assign mesh_7_7_io_in_valid_0 = _T_511_0; // @[Mesh.scala 78:26:example.TestHarness.GemminiSocTest1RocketConfig864.fir@180142.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_0 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1_0 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2_0 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3_0 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_4_0 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_5_0 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_6_0 = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_7_0 = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_8_0 = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_9_0 = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_10_0 = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_11_0 = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_12_0 = _RAND_12[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_13_0 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_14_0 = _RAND_14[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_15_0 = _RAND_15[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_16_0 = _RAND_16[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_17_0 = _RAND_17[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_18_0 = _RAND_18[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_19_0 = _RAND_19[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_20_0 = _RAND_20[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_21_0 = _RAND_21[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_22_0 = _RAND_22[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_23_0 = _RAND_23[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_24_0 = _RAND_24[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_25_0 = _RAND_25[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_26_0 = _RAND_26[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_27_0 = _RAND_27[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_28_0 = _RAND_28[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_29_0 = _RAND_29[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_30_0 = _RAND_30[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_31_0 = _RAND_31[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_32_0 = _RAND_32[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_33_0 = _RAND_33[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_34_0 = _RAND_34[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_35_0 = _RAND_35[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_36_0 = _RAND_36[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_37_0 = _RAND_37[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_38_0 = _RAND_38[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_39_0 = _RAND_39[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_40_0 = _RAND_40[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_41_0 = _RAND_41[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_42_0 = _RAND_42[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_43_0 = _RAND_43[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_44_0 = _RAND_44[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_45_0 = _RAND_45[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_46_0 = _RAND_46[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_47_0 = _RAND_47[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_48_0 = _RAND_48[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_49_0 = _RAND_49[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_50_0 = _RAND_50[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_51_0 = _RAND_51[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_52_0 = _RAND_52[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_53_0 = _RAND_53[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_54_0 = _RAND_54[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_55_0 = _RAND_55[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_56_0 = _RAND_56[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_57_0 = _RAND_57[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_58_0 = _RAND_58[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_59_0 = _RAND_59[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_60_0 = _RAND_60[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_61_0 = _RAND_61[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_62_0 = _RAND_62[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_63_0 = _RAND_63[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_64_0 = _RAND_64[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_65_0 = _RAND_65[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_66_0 = _RAND_66[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_67_0 = _RAND_67[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_68_0 = _RAND_68[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_69_0 = _RAND_69[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_70_0 = _RAND_70[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_71_0 = _RAND_71[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_72_0 = _RAND_72[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_73_0 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_74_0 = _RAND_74[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_75_0 = _RAND_75[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_76_0 = _RAND_76[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_77_0 = _RAND_77[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_78_0 = _RAND_78[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_79_0 = _RAND_79[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_80_0 = _RAND_80[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_81_0 = _RAND_81[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_82_0 = _RAND_82[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_83_0 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_84_0 = _RAND_84[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_85_0 = _RAND_85[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_86_0 = _RAND_86[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_87_0 = _RAND_87[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_88_0 = _RAND_88[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_89_0 = _RAND_89[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_90_0 = _RAND_90[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_91_0 = _RAND_91[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_92_0 = _RAND_92[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_93_0 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_94_0 = _RAND_94[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_95_0 = _RAND_95[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_96_0 = _RAND_96[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_97_0 = _RAND_97[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_98_0 = _RAND_98[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_99_0 = _RAND_99[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_100_0 = _RAND_100[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_101_0 = _RAND_101[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_102_0 = _RAND_102[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_103_0 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_104_0 = _RAND_104[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_105_0 = _RAND_105[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_106_0 = _RAND_106[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_107_0 = _RAND_107[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_108_0 = _RAND_108[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_109_0 = _RAND_109[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_110_0 = _RAND_110[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_111_0 = _RAND_111[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_112_0 = _RAND_112[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_113_0 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_114_0 = _RAND_114[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_115_0 = _RAND_115[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_116_0 = _RAND_116[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_117_0 = _RAND_117[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_118_0 = _RAND_118[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_119_0 = _RAND_119[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_120_0 = _RAND_120[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_121_0 = _RAND_121[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_122_0 = _RAND_122[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_123_0 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_124_0 = _RAND_124[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_125_0 = _RAND_125[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_126_0 = _RAND_126[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_127_0 = _RAND_127[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_128_0 = _RAND_128[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_129_0 = _RAND_129[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_130_0 = _RAND_130[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_131_0 = _RAND_131[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_132_0 = _RAND_132[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_133_0 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_134_0 = _RAND_134[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_135_0 = _RAND_135[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_136_0 = _RAND_136[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_137_0 = _RAND_137[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_138_0 = _RAND_138[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_139_0 = _RAND_139[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_140_0 = _RAND_140[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_141_0 = _RAND_141[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_142_0 = _RAND_142[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_143_0 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_144_0 = _RAND_144[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_145_0 = _RAND_145[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_146_0 = _RAND_146[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_147_0 = _RAND_147[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_148_0 = _RAND_148[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_149_0 = _RAND_149[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_150_0 = _RAND_150[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_151_0 = _RAND_151[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_152_0 = _RAND_152[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_153_0 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_154_0 = _RAND_154[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_155_0 = _RAND_155[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_156_0 = _RAND_156[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_157_0 = _RAND_157[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_158_0 = _RAND_158[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_159_0 = _RAND_159[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_160_0 = _RAND_160[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_161_0 = _RAND_161[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_162_0 = _RAND_162[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_163_0 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_164_0 = _RAND_164[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_165_0 = _RAND_165[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_166_0 = _RAND_166[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_167_0 = _RAND_167[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_168_0 = _RAND_168[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_169_0 = _RAND_169[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_170_0 = _RAND_170[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_171_0 = _RAND_171[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_172_0 = _RAND_172[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_173_0 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_174_0 = _RAND_174[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_175_0 = _RAND_175[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_176_0 = _RAND_176[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_177_0 = _RAND_177[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_178_0 = _RAND_178[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_179_0 = _RAND_179[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_180_0 = _RAND_180[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_181_0 = _RAND_181[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_182_0 = _RAND_182[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_183_0 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_184_0 = _RAND_184[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_185_0 = _RAND_185[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_186_0 = _RAND_186[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_187_0 = _RAND_187[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_188_0 = _RAND_188[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_189_0 = _RAND_189[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_190_0 = _RAND_190[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_191_0 = _RAND_191[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_192_0 = _RAND_192[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_193_0 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_194_0 = _RAND_194[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_195_0 = _RAND_195[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_196_0 = _RAND_196[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_197_0 = _RAND_197[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_198_0 = _RAND_198[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_199_0 = _RAND_199[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_200_0 = _RAND_200[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_201_0 = _RAND_201[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_202_0 = _RAND_202[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_203_0 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_204_0 = _RAND_204[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_205_0 = _RAND_205[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_206_0 = _RAND_206[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_207_0 = _RAND_207[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_208_0 = _RAND_208[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_209_0 = _RAND_209[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_210_0 = _RAND_210[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_211_0 = _RAND_211[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_212_0 = _RAND_212[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_213_0 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_214_0 = _RAND_214[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_215_0 = _RAND_215[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_216_0 = _RAND_216[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_217_0 = _RAND_217[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_218_0 = _RAND_218[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_219_0 = _RAND_219[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_220_0 = _RAND_220[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_221_0 = _RAND_221[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_222_0 = _RAND_222[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_223_0 = _RAND_223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_224_0 = _RAND_224[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_225_0 = _RAND_225[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_226_0 = _RAND_226[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_227_0 = _RAND_227[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_228_0 = _RAND_228[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_229_0 = _RAND_229[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_230_0 = _RAND_230[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_231_0 = _RAND_231[(dbits-1):0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_232_0_propagate = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_232_0_shift = _RAND_233[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_233_0 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_234 = _RAND_235[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_236 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_237 = _RAND_237[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_239 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_240 = _RAND_239[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_242 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_243 = _RAND_241[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_245 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_246 = _RAND_243[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_248 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_249 = _RAND_245[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_251 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_252 = _RAND_247[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_254 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_255 = _RAND_249[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_257 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_258_0_propagate = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_258_0_shift = _RAND_252[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_259_0 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_260 = _RAND_254[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_262 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_263 = _RAND_256[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_265 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_266 = _RAND_258[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_268 = _RAND_259[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_269 = _RAND_260[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_271 = _RAND_261[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _T_272 = _RAND_262[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _T_274 = _RAND_263[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _T_275 = _RAND_264[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _T_277 = _RAND_265[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _T_278 = _RAND_266[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _T_280 = _RAND_267[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _T_281 = _RAND_268[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _T_283 = _RAND_269[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _T_284_0_propagate = _RAND_270[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_284_0_shift = _RAND_271[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_285_0 = _RAND_272[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _T_286 = _RAND_273[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_288 = _RAND_274[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _T_289 = _RAND_275[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_291 = _RAND_276[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_292 = _RAND_277[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_294 = _RAND_278[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _T_295 = _RAND_279[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_297 = _RAND_280[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _T_298 = _RAND_281[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _T_300 = _RAND_282[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_301 = _RAND_283[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_303 = _RAND_284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _T_304 = _RAND_285[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _T_306 = _RAND_286[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _T_307 = _RAND_287[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _T_309 = _RAND_288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _T_310_0_propagate = _RAND_289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _T_310_0_shift = _RAND_290[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _T_311_0 = _RAND_291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _T_312 = _RAND_292[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _T_314 = _RAND_293[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _T_315 = _RAND_294[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _T_317 = _RAND_295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _T_318 = _RAND_296[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _T_320 = _RAND_297[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _T_321 = _RAND_298[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _T_323 = _RAND_299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _T_324 = _RAND_300[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _T_326 = _RAND_301[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _T_327 = _RAND_302[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _T_329 = _RAND_303[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _T_330 = _RAND_304[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _T_332 = _RAND_305[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _T_333 = _RAND_306[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _T_335 = _RAND_307[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _T_336_0_propagate = _RAND_308[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _T_336_0_shift = _RAND_309[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _T_337_0 = _RAND_310[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _T_338 = _RAND_311[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _T_340 = _RAND_312[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _T_341 = _RAND_313[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _T_343 = _RAND_314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _T_344 = _RAND_315[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _T_346 = _RAND_316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _T_347 = _RAND_317[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _T_349 = _RAND_318[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _T_350 = _RAND_319[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _T_352 = _RAND_320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _T_353 = _RAND_321[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _T_355 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _T_356 = _RAND_323[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _T_358 = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _T_359 = _RAND_325[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _T_361 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _T_362_0_propagate = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _T_362_0_shift = _RAND_328[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _T_363_0 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _T_364 = _RAND_330[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _T_366 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _T_367 = _RAND_332[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _T_369 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _T_370 = _RAND_334[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _T_372 = _RAND_335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _T_373 = _RAND_336[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _T_375 = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _T_376 = _RAND_338[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _T_378 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _T_379 = _RAND_340[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _T_381 = _RAND_341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _T_382 = _RAND_342[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _T_384 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _T_385 = _RAND_344[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _T_387 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _T_388_0_propagate = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _T_388_0_shift = _RAND_347[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _T_389_0 = _RAND_348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _T_390 = _RAND_349[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _T_392 = _RAND_350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _T_393 = _RAND_351[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _T_395 = _RAND_352[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _T_396 = _RAND_353[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _T_398 = _RAND_354[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _T_399 = _RAND_355[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _T_401 = _RAND_356[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _T_402 = _RAND_357[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _T_404 = _RAND_358[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _T_405 = _RAND_359[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _T_407 = _RAND_360[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _T_408 = _RAND_361[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _T_410 = _RAND_362[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _T_411 = _RAND_363[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _T_413 = _RAND_364[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _T_414_0_propagate = _RAND_365[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _T_414_0_shift = _RAND_366[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _T_415_0 = _RAND_367[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _T_416 = _RAND_368[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _T_418 = _RAND_369[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _T_419 = _RAND_370[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _T_421 = _RAND_371[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _T_422 = _RAND_372[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _T_424 = _RAND_373[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _T_425 = _RAND_374[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _T_427 = _RAND_375[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _T_428 = _RAND_376[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _T_430 = _RAND_377[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _T_431 = _RAND_378[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  _T_433 = _RAND_379[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  _T_434 = _RAND_380[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _T_436 = _RAND_381[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  _T_437 = _RAND_382[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  _T_439 = _RAND_383[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  _T_440_0 = _RAND_384[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  _T_441_0 = _RAND_385[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  _T_442_0 = _RAND_386[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  _T_443_0 = _RAND_387[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  _T_444_0 = _RAND_388[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  _T_445_0 = _RAND_389[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  _T_446_0 = _RAND_390[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  _T_447_0 = _RAND_391[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  _T_448_0 = _RAND_392[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  _T_449_0 = _RAND_393[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  _T_450_0 = _RAND_394[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  _T_451_0 = _RAND_395[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  _T_452_0 = _RAND_396[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  _T_453_0 = _RAND_397[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  _T_454_0 = _RAND_398[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  _T_455_0 = _RAND_399[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  _T_456_0 = _RAND_400[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  _T_457_0 = _RAND_401[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  _T_458_0 = _RAND_402[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  _T_459_0 = _RAND_403[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  _T_460_0 = _RAND_404[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  _T_461_0 = _RAND_405[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  _T_462_0 = _RAND_406[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  _T_463_0 = _RAND_407[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  _T_464_0 = _RAND_408[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  _T_465_0 = _RAND_409[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  _T_466_0 = _RAND_410[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  _T_467_0 = _RAND_411[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  _T_468_0 = _RAND_412[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  _T_469_0 = _RAND_413[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  _T_470_0 = _RAND_414[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  _T_471_0 = _RAND_415[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  _T_472_0 = _RAND_416[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  _T_473_0 = _RAND_417[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  _T_474_0 = _RAND_418[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  _T_475_0 = _RAND_419[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  _T_476_0 = _RAND_420[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  _T_477_0 = _RAND_421[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  _T_478_0 = _RAND_422[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  _T_479_0 = _RAND_423[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  _T_480_0 = _RAND_424[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  _T_481_0 = _RAND_425[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  _T_482_0 = _RAND_426[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  _T_483_0 = _RAND_427[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  _T_484_0 = _RAND_428[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  _T_485_0 = _RAND_429[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  _T_486_0 = _RAND_430[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  _T_487_0 = _RAND_431[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  _T_488_0 = _RAND_432[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  _T_489_0 = _RAND_433[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  _T_490_0 = _RAND_434[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  _T_491_0 = _RAND_435[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  _T_492_0 = _RAND_436[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  _T_493_0 = _RAND_437[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  _T_494_0 = _RAND_438[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  _T_495_0 = _RAND_439[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  _T_496_0 = _RAND_440[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  _T_497_0 = _RAND_441[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  _T_498_0 = _RAND_442[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  _T_499_0 = _RAND_443[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  _T_500_0 = _RAND_444[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  _T_501_0 = _RAND_445[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  _T_502_0 = _RAND_446[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  _T_503_0 = _RAND_447[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  _T_504_0 = _RAND_448[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  _T_505_0 = _RAND_449[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  _T_506_0 = _RAND_450[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  _T_507_0 = _RAND_451[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  _T_508_0 = _RAND_452[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  _T_509_0 = _RAND_453[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  _T_510_0 = _RAND_454[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  _T_511_0 = _RAND_455[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    //_T_0 <= io_in_a_0_0;
    _T_1_0 <= io_in_a_0_0;
    _T_2_0 <= mesh_0_0_io_out_a_0;
    _T_3_0 <= mesh_0_1_io_out_a_0;
    _T_4_0 <= mesh_0_2_io_out_a_0;
    _T_5_0 <= mesh_0_3_io_out_a_0;
    _T_6_0 <= mesh_0_4_io_out_a_0;
    _T_7_0 <= mesh_0_5_io_out_a_0;
    _T_8_0 <= mesh_0_6_io_out_a_0;
    //_T_9_0 <= io_in_a_1_0;
    _T_10_0 <= io_in_a_1_0;
    _T_11_0 <= mesh_1_0_io_out_a_0;
    _T_12_0 <= mesh_1_1_io_out_a_0;
    _T_13_0 <= mesh_1_2_io_out_a_0;
    _T_14_0 <= mesh_1_3_io_out_a_0;
    _T_15_0 <= mesh_1_4_io_out_a_0;
    _T_16_0 <= mesh_1_5_io_out_a_0;
    _T_17_0 <= mesh_1_6_io_out_a_0;
    //_T_18_0 <= io_in_a_2_0;
    _T_19_0 <= io_in_a_2_0;
    _T_20_0 <= mesh_2_0_io_out_a_0;
    _T_21_0 <= mesh_2_1_io_out_a_0;
    _T_22_0 <= mesh_2_2_io_out_a_0;
    _T_23_0 <= mesh_2_3_io_out_a_0;
    _T_24_0 <= mesh_2_4_io_out_a_0;
    _T_25_0 <= mesh_2_5_io_out_a_0;
    _T_26_0 <= mesh_2_6_io_out_a_0;
    //_T_27_0 <= io_in_a_3_0;
    _T_28_0 <= io_in_a_3_0;
    _T_29_0 <= mesh_3_0_io_out_a_0;
    _T_30_0 <= mesh_3_1_io_out_a_0;
    _T_31_0 <= mesh_3_2_io_out_a_0;
    _T_32_0 <= mesh_3_3_io_out_a_0;
    _T_33_0 <= mesh_3_4_io_out_a_0;
    _T_34_0 <= mesh_3_5_io_out_a_0;
    _T_35_0 <= mesh_3_6_io_out_a_0;
    //_T_36_0 <= io_in_a_4_0;
    _T_37_0 <= io_in_a_4_0;
    _T_38_0 <= mesh_4_0_io_out_a_0;
    _T_39_0 <= mesh_4_1_io_out_a_0;
    _T_40_0 <= mesh_4_2_io_out_a_0;
    _T_41_0 <= mesh_4_3_io_out_a_0;
    _T_42_0 <= mesh_4_4_io_out_a_0;
    _T_43_0 <= mesh_4_5_io_out_a_0;
    _T_44_0 <= mesh_4_6_io_out_a_0;
    //_T_45_0 <= io_in_a_5_0;
    _T_46_0 <= io_in_a_5_0;
    _T_47_0 <= mesh_5_0_io_out_a_0;
    _T_48_0 <= mesh_5_1_io_out_a_0;
    _T_49_0 <= mesh_5_2_io_out_a_0;
    _T_50_0 <= mesh_5_3_io_out_a_0;
    _T_51_0 <= mesh_5_4_io_out_a_0;
    _T_52_0 <= mesh_5_5_io_out_a_0;
    _T_53_0 <= mesh_5_6_io_out_a_0;
    //_T_54_0 <= io_in_a_6_0;
    _T_55_0 <= io_in_a_6_0;
    _T_56_0 <= mesh_6_0_io_out_a_0;
    _T_57_0 <= mesh_6_1_io_out_a_0;
    _T_58_0 <= mesh_6_2_io_out_a_0;
    _T_59_0 <= mesh_6_3_io_out_a_0;
    _T_60_0 <= mesh_6_4_io_out_a_0;
    _T_61_0 <= mesh_6_5_io_out_a_0;
    _T_62_0 <= mesh_6_6_io_out_a_0;
    //_T_63_0 <= io_in_a_7_0;
    _T_64_0 <= io_in_a_7_0;
    _T_65_0 <= mesh_7_0_io_out_a_0;
    _T_66_0 <= mesh_7_1_io_out_a_0;
    _T_67_0 <= mesh_7_2_io_out_a_0;
    _T_68_0 <= mesh_7_3_io_out_a_0;
    _T_69_0 <= mesh_7_4_io_out_a_0;
    _T_70_0 <= mesh_7_5_io_out_a_0;
    _T_71_0 <= mesh_7_6_io_out_a_0;
    //_T_72_0 <= io_in_d_0_0;
    //_T_73_0 <= io_in_valid_0_0;
     if (io_in_valid_0_0) begin
    _T_74_0 <= io_in_d_0_0;
    end
    if (mesh_0_0_io_out_valid_0) begin
      _T_75_0 <= mesh_0_0_io_out_b_0;
    end
    if (mesh_1_0_io_out_valid_0) begin
      _T_76_0 <= mesh_1_0_io_out_b_0;
    end
    if (mesh_2_0_io_out_valid_0) begin
      _T_77_0 <= mesh_2_0_io_out_b_0;
    end
    if (mesh_3_0_io_out_valid_0) begin
      _T_78_0 <= mesh_3_0_io_out_b_0;
    end
    if (mesh_4_0_io_out_valid_0) begin
      _T_79_0 <= mesh_4_0_io_out_b_0;
    end
    if (mesh_5_0_io_out_valid_0) begin
      _T_80_0 <= mesh_5_0_io_out_b_0;
    end
    if (mesh_6_0_io_out_valid_0) begin
      _T_81_0 <= mesh_6_0_io_out_b_0;
    end
    //_T_82_0 <= io_in_d_1_0;
    //_T_83_0 <= io_in_valid_1_0;
     if (io_in_valid_1_0) begin
    _T_84_0 <= io_in_d_1_0;
    end
    if (mesh_0_1_io_out_valid_0) begin
      _T_85_0 <= mesh_0_1_io_out_b_0;
    end
    if (mesh_1_1_io_out_valid_0) begin
      _T_86_0 <= mesh_1_1_io_out_b_0;
    end
    if (mesh_2_1_io_out_valid_0) begin
      _T_87_0 <= mesh_2_1_io_out_b_0;
    end
    if (mesh_3_1_io_out_valid_0) begin
      _T_88_0 <= mesh_3_1_io_out_b_0;
    end
    if (mesh_4_1_io_out_valid_0) begin
      _T_89_0 <= mesh_4_1_io_out_b_0;
    end
    if (mesh_5_1_io_out_valid_0) begin
      _T_90_0 <= mesh_5_1_io_out_b_0;
    end
    if (mesh_6_1_io_out_valid_0) begin
      _T_91_0 <= mesh_6_1_io_out_b_0;
    end
    //_T_92_0 <= io_in_d_2_0;
    //_T_93_0 <= io_in_valid_2_0;
     if (io_in_valid_2_0) begin
    _T_94_0 <= io_in_d_2_0;
    end
    if (mesh_0_2_io_out_valid_0) begin
      _T_95_0 <= mesh_0_2_io_out_b_0;
    end
    if (mesh_1_2_io_out_valid_0) begin
      _T_96_0 <= mesh_1_2_io_out_b_0;
    end
    if (mesh_2_2_io_out_valid_0) begin
      _T_97_0 <= mesh_2_2_io_out_b_0;
    end
    if (mesh_3_2_io_out_valid_0) begin
      _T_98_0 <= mesh_3_2_io_out_b_0;
    end
    if (mesh_4_2_io_out_valid_0) begin
      _T_99_0 <= mesh_4_2_io_out_b_0;
    end
    if (mesh_5_2_io_out_valid_0) begin
      _T_100_0 <= mesh_5_2_io_out_b_0;
    end
    if (mesh_6_2_io_out_valid_0) begin
      _T_101_0 <= mesh_6_2_io_out_b_0;
    end
    //_T_102_0 <= io_in_d_3_0;
    //_T_103_0 <= io_in_valid_3_0;
     if (io_in_valid_3_0) begin
    _T_104_0 <= io_in_d_3_0;
    end
    if (mesh_0_3_io_out_valid_0) begin
      _T_105_0 <= mesh_0_3_io_out_b_0;
    end
    if (mesh_1_3_io_out_valid_0) begin
      _T_106_0 <= mesh_1_3_io_out_b_0;
    end
    if (mesh_2_3_io_out_valid_0) begin
      _T_107_0 <= mesh_2_3_io_out_b_0;
    end
    if (mesh_3_3_io_out_valid_0) begin
      _T_108_0 <= mesh_3_3_io_out_b_0;
    end
    if (mesh_4_3_io_out_valid_0) begin
      _T_109_0 <= mesh_4_3_io_out_b_0;
    end
    if (mesh_5_3_io_out_valid_0) begin
      _T_110_0 <= mesh_5_3_io_out_b_0;
    end
    if (mesh_6_3_io_out_valid_0) begin
      _T_111_0 <= mesh_6_3_io_out_b_0;
    end
    //_T_112_0 <= io_in_d_4_0;
    //_T_113_0 <= io_in_valid_4_0;
     if (io_in_valid_4_0) begin
    _T_114_0 <= io_in_d_4_0;
    end
    if (mesh_0_4_io_out_valid_0) begin
      _T_115_0 <= mesh_0_4_io_out_b_0;
    end
    if (mesh_1_4_io_out_valid_0) begin
      _T_116_0 <= mesh_1_4_io_out_b_0;
    end
    if (mesh_2_4_io_out_valid_0) begin
      _T_117_0 <= mesh_2_4_io_out_b_0;
    end
    if (mesh_3_4_io_out_valid_0) begin
      _T_118_0 <= mesh_3_4_io_out_b_0;
    end
    if (mesh_4_4_io_out_valid_0) begin
      _T_119_0 <= mesh_4_4_io_out_b_0;
    end
    if (mesh_5_4_io_out_valid_0) begin
      _T_120_0 <= mesh_5_4_io_out_b_0;
    end
    if (mesh_6_4_io_out_valid_0) begin
      _T_121_0 <= mesh_6_4_io_out_b_0;
    end
    //_T_122_0 <= io_in_d_5_0;
    //_T_123_0 <= io_in_valid_5_0;
     if (io_in_valid_5_0) begin
    _T_124_0 <= io_in_d_5_0;
    end
    if (mesh_0_5_io_out_valid_0) begin
      _T_125_0 <= mesh_0_5_io_out_b_0;
    end
    if (mesh_1_5_io_out_valid_0) begin
      _T_126_0 <= mesh_1_5_io_out_b_0;
    end
    if (mesh_2_5_io_out_valid_0) begin
      _T_127_0 <= mesh_2_5_io_out_b_0;
    end
    if (mesh_3_5_io_out_valid_0) begin
      _T_128_0 <= mesh_3_5_io_out_b_0;
    end
    if (mesh_4_5_io_out_valid_0) begin
      _T_129_0 <= mesh_4_5_io_out_b_0;
    end
    if (mesh_5_5_io_out_valid_0) begin
      _T_130_0 <= mesh_5_5_io_out_b_0;
    end
    if (mesh_6_5_io_out_valid_0) begin
      _T_131_0 <= mesh_6_5_io_out_b_0;
    end
    //_T_132_0 <= io_in_d_6_0;
    //_T_133_0 <= io_in_valid_6_0;
     if (io_in_valid_6_0) begin
    _T_134_0 <= io_in_d_6_0;
    end
    if (mesh_0_6_io_out_valid_0) begin
      _T_135_0 <= mesh_0_6_io_out_b_0;
    end
    if (mesh_1_6_io_out_valid_0) begin
      _T_136_0 <= mesh_1_6_io_out_b_0;
    end
    if (mesh_2_6_io_out_valid_0) begin
      _T_137_0 <= mesh_2_6_io_out_b_0;
    end
    if (mesh_3_6_io_out_valid_0) begin
      _T_138_0 <= mesh_3_6_io_out_b_0;
    end
    if (mesh_4_6_io_out_valid_0) begin
      _T_139_0 <= mesh_4_6_io_out_b_0;
    end
    if (mesh_5_6_io_out_valid_0) begin
      _T_140_0 <= mesh_5_6_io_out_b_0;
    end
    if (mesh_6_6_io_out_valid_0) begin
      _T_141_0 <= mesh_6_6_io_out_b_0;
    end
    //_T_142_0 <= io_in_d_7_0;
    //_T_143_0 <= io_in_valid_7_0;
     if (io_in_valid_7_0) begin
    _T_144_0 <= io_in_d_7_0;
    end
    if (mesh_0_7_io_out_valid_0) begin
      _T_145_0 <= mesh_0_7_io_out_b_0;
    end
    if (mesh_1_7_io_out_valid_0) begin
      _T_146_0 <= mesh_1_7_io_out_b_0;
    end
    if (mesh_2_7_io_out_valid_0) begin
      _T_147_0 <= mesh_2_7_io_out_b_0;
    end
    if (mesh_3_7_io_out_valid_0) begin
      _T_148_0 <= mesh_3_7_io_out_b_0;
    end
    if (mesh_4_7_io_out_valid_0) begin
      _T_149_0 <= mesh_4_7_io_out_b_0;
    end
    if (mesh_5_7_io_out_valid_0) begin
      _T_150_0 <= mesh_5_7_io_out_b_0;
    end
    if (mesh_6_7_io_out_valid_0) begin
      _T_151_0 <= mesh_6_7_io_out_b_0;
    end
    //_T_152_0 <= io_in_b_0_0;
    //_T_153_0 <= io_in_valid_0_0;
     if (io_in_valid_0_0) begin
    _T_154_0 <= io_in_b_0_0;
    end
    if (mesh_0_0_io_out_valid_0) begin
      _T_155_0 <= mesh_0_0_io_out_c_0;
    end
    if (mesh_1_0_io_out_valid_0) begin
      _T_156_0 <= mesh_1_0_io_out_c_0;
    end
    if (mesh_2_0_io_out_valid_0) begin
      _T_157_0 <= mesh_2_0_io_out_c_0;
    end
    if (mesh_3_0_io_out_valid_0) begin
      _T_158_0 <= mesh_3_0_io_out_c_0;
    end
    if (mesh_4_0_io_out_valid_0) begin
      _T_159_0 <= mesh_4_0_io_out_c_0;
    end
    if (mesh_5_0_io_out_valid_0) begin
      _T_160_0 <= mesh_5_0_io_out_c_0;
    end
    if (mesh_6_0_io_out_valid_0) begin
      _T_161_0 <= mesh_6_0_io_out_c_0;
    end
    //_T_162_0 <= io_in_b_1_0;
    //_T_163_0 <= io_in_valid_1_0;
     if (io_in_valid_1_0) begin
    _T_164_0 <= io_in_b_1_0;
    end
    if (mesh_0_1_io_out_valid_0) begin
      _T_165_0 <= mesh_0_1_io_out_c_0;
    end
    if (mesh_1_1_io_out_valid_0) begin
      _T_166_0 <= mesh_1_1_io_out_c_0;
    end
    if (mesh_2_1_io_out_valid_0) begin
      _T_167_0 <= mesh_2_1_io_out_c_0;
    end
    if (mesh_3_1_io_out_valid_0) begin
      _T_168_0 <= mesh_3_1_io_out_c_0;
    end
    if (mesh_4_1_io_out_valid_0) begin
      _T_169_0 <= mesh_4_1_io_out_c_0;
    end
    if (mesh_5_1_io_out_valid_0) begin
      _T_170_0 <= mesh_5_1_io_out_c_0;
    end
    if (mesh_6_1_io_out_valid_0) begin
      _T_171_0 <= mesh_6_1_io_out_c_0;
    end
    //_T_172_0 <= io_in_b_2_0;
    //_T_173_0 <= io_in_valid_2_0;
     if (io_in_valid_2_0) begin
    _T_174_0 <= io_in_b_2_0;
    end
    if (mesh_0_2_io_out_valid_0) begin
      _T_175_0 <= mesh_0_2_io_out_c_0;
    end
    if (mesh_1_2_io_out_valid_0) begin
      _T_176_0 <= mesh_1_2_io_out_c_0;
    end
    if (mesh_2_2_io_out_valid_0) begin
      _T_177_0 <= mesh_2_2_io_out_c_0;
    end
    if (mesh_3_2_io_out_valid_0) begin
      _T_178_0 <= mesh_3_2_io_out_c_0;
    end
    if (mesh_4_2_io_out_valid_0) begin
      _T_179_0 <= mesh_4_2_io_out_c_0;
    end
    if (mesh_5_2_io_out_valid_0) begin
      _T_180_0 <= mesh_5_2_io_out_c_0;
    end
    if (mesh_6_2_io_out_valid_0) begin
      _T_181_0 <= mesh_6_2_io_out_c_0;
    end
    //_T_182_0 <= io_in_b_3_0;
    //_T_183_0 <= io_in_valid_3_0;
     if (io_in_valid_3_0) begin
    _T_184_0 <= io_in_b_3_0;
    end
    if (mesh_0_3_io_out_valid_0) begin
      _T_185_0 <= mesh_0_3_io_out_c_0;
    end
    if (mesh_1_3_io_out_valid_0) begin
      _T_186_0 <= mesh_1_3_io_out_c_0;
    end
    if (mesh_2_3_io_out_valid_0) begin
      _T_187_0 <= mesh_2_3_io_out_c_0;
    end
    if (mesh_3_3_io_out_valid_0) begin
      _T_188_0 <= mesh_3_3_io_out_c_0;
    end
    if (mesh_4_3_io_out_valid_0) begin
      _T_189_0 <= mesh_4_3_io_out_c_0;
    end
    if (mesh_5_3_io_out_valid_0) begin
      _T_190_0 <= mesh_5_3_io_out_c_0;
    end
    if (mesh_6_3_io_out_valid_0) begin
      _T_191_0 <= mesh_6_3_io_out_c_0;
    end
    //_T_192_0 <= io_in_b_4_0;
    //_T_193_0 <= io_in_valid_4_0;
     if (io_in_valid_4_0) begin
    _T_194_0 <= io_in_b_4_0;
    end
    if (mesh_0_4_io_out_valid_0) begin
      _T_195_0 <= mesh_0_4_io_out_c_0;
    end
    if (mesh_1_4_io_out_valid_0) begin
      _T_196_0 <= mesh_1_4_io_out_c_0;
    end
    if (mesh_2_4_io_out_valid_0) begin
      _T_197_0 <= mesh_2_4_io_out_c_0;
    end
    if (mesh_3_4_io_out_valid_0) begin
      _T_198_0 <= mesh_3_4_io_out_c_0;
    end
    if (mesh_4_4_io_out_valid_0) begin
      _T_199_0 <= mesh_4_4_io_out_c_0;
    end
    if (mesh_5_4_io_out_valid_0) begin
      _T_200_0 <= mesh_5_4_io_out_c_0;
    end
    if (mesh_6_4_io_out_valid_0) begin
      _T_201_0 <= mesh_6_4_io_out_c_0;
    end
    //_T_202_0 <= io_in_b_5_0;
    //_T_203_0 <= io_in_valid_5_0;
     if (io_in_valid_5_0) begin
    _T_204_0 <= io_in_b_5_0;
    end
    if (mesh_0_5_io_out_valid_0) begin
      _T_205_0 <= mesh_0_5_io_out_c_0;
    end
    if (mesh_1_5_io_out_valid_0) begin
      _T_206_0 <= mesh_1_5_io_out_c_0;
    end
    if (mesh_2_5_io_out_valid_0) begin
      _T_207_0 <= mesh_2_5_io_out_c_0;
    end
    if (mesh_3_5_io_out_valid_0) begin
      _T_208_0 <= mesh_3_5_io_out_c_0;
    end
    if (mesh_4_5_io_out_valid_0) begin
      _T_209_0 <= mesh_4_5_io_out_c_0;
    end
    if (mesh_5_5_io_out_valid_0) begin
      _T_210_0 <= mesh_5_5_io_out_c_0;
    end
    if (mesh_6_5_io_out_valid_0) begin
      _T_211_0 <= mesh_6_5_io_out_c_0;
    end
    //_T_212_0 <= io_in_b_6_0;
    //_T_213_0 <= io_in_valid_6_0;
     if (io_in_valid_6_0) begin
    _T_214_0 <= io_in_b_6_0;
    end
    if (mesh_0_6_io_out_valid_0) begin
      _T_215_0 <= mesh_0_6_io_out_c_0;
    end
    if (mesh_1_6_io_out_valid_0) begin
      _T_216_0 <= mesh_1_6_io_out_c_0;
    end
    if (mesh_2_6_io_out_valid_0) begin
      _T_217_0 <= mesh_2_6_io_out_c_0;
    end
    if (mesh_3_6_io_out_valid_0) begin
      _T_218_0 <= mesh_3_6_io_out_c_0;
    end
    if (mesh_4_6_io_out_valid_0) begin
      _T_219_0 <= mesh_4_6_io_out_c_0;
    end
    if (mesh_5_6_io_out_valid_0) begin
      _T_220_0 <= mesh_5_6_io_out_c_0;
    end
    if (mesh_6_6_io_out_valid_0) begin
      _T_221_0 <= mesh_6_6_io_out_c_0;
    end
    //_T_222_0 <= io_in_b_7_0;
    //_T_223_0 <= io_in_valid_7_0;
     if (io_in_valid_7_0) begin
    _T_224_0 <= io_in_b_7_0;
    end
    if (mesh_0_7_io_out_valid_0) begin
      _T_225_0 <= mesh_0_7_io_out_c_0;
    end
    if (mesh_1_7_io_out_valid_0) begin
      _T_226_0 <= mesh_1_7_io_out_c_0;
    end
    if (mesh_2_7_io_out_valid_0) begin
      _T_227_0 <= mesh_2_7_io_out_c_0;
    end
    if (mesh_3_7_io_out_valid_0) begin
      _T_228_0 <= mesh_3_7_io_out_c_0;
    end
    if (mesh_4_7_io_out_valid_0) begin
      _T_229_0 <= mesh_4_7_io_out_c_0;
    end
    if (mesh_5_7_io_out_valid_0) begin
      _T_230_0 <= mesh_5_7_io_out_c_0;
    end
    if (mesh_6_7_io_out_valid_0) begin
      _T_231_0 <= mesh_6_7_io_out_c_0;
    end
    //_T_232_0_propagate <= io_in_control_0_0_propagate;
    //_T_232_0_shift <= io_in_control_0_0_shift;
    //_T_233_0 <= io_in_valid_0_0;
     if (io_in_valid_0_0) begin
    _T_234 <= io_in_control_0_0_shift;
    end
     if (io_in_valid_0_0) begin
    _T_236 <= io_in_control_0_0_propagate;
    end
    if (mesh_0_0_io_out_valid_0) begin
      _T_237 <= mesh_0_0_io_out_control_0_shift;
    end
    if (mesh_0_0_io_out_valid_0) begin
      _T_239 <= mesh_0_0_io_out_control_0_propagate;
    end
    if (mesh_1_0_io_out_valid_0) begin
      _T_240 <= mesh_1_0_io_out_control_0_shift;
    end
    if (mesh_1_0_io_out_valid_0) begin
      _T_242 <= mesh_1_0_io_out_control_0_propagate;
    end
    if (mesh_2_0_io_out_valid_0) begin
      _T_243 <= mesh_2_0_io_out_control_0_shift;
    end
    if (mesh_2_0_io_out_valid_0) begin
      _T_245 <= mesh_2_0_io_out_control_0_propagate;
    end
    if (mesh_3_0_io_out_valid_0) begin
      _T_246 <= mesh_3_0_io_out_control_0_shift;
    end
    if (mesh_3_0_io_out_valid_0) begin
      _T_248 <= mesh_3_0_io_out_control_0_propagate;
    end
    if (mesh_4_0_io_out_valid_0) begin
      _T_249 <= mesh_4_0_io_out_control_0_shift;
    end
    if (mesh_4_0_io_out_valid_0) begin
      _T_251 <= mesh_4_0_io_out_control_0_propagate;
    end
    if (mesh_5_0_io_out_valid_0) begin
      _T_252 <= mesh_5_0_io_out_control_0_shift;
    end
    if (mesh_5_0_io_out_valid_0) begin
      _T_254 <= mesh_5_0_io_out_control_0_propagate;
    end
    if (mesh_6_0_io_out_valid_0) begin
      _T_255 <= mesh_6_0_io_out_control_0_shift;
    end
    if (mesh_6_0_io_out_valid_0) begin
      _T_257 <= mesh_6_0_io_out_control_0_propagate;
    end
    //_T_258_0_propagate <= io_in_control_1_0_propagate;
    //_T_258_0_shift <= io_in_control_1_0_shift;
    //_T_259_0 <= io_in_valid_1_0;
     if (io_in_valid_1_0) begin
    _T_260 <= io_in_control_1_0_shift;
    end
     if (io_in_valid_1_0) begin
    _T_262 <= io_in_control_1_0_propagate;
    end
    if (mesh_0_1_io_out_valid_0) begin
      _T_263 <= mesh_0_1_io_out_control_0_shift;
    end
    if (mesh_0_1_io_out_valid_0) begin
      _T_265 <= mesh_0_1_io_out_control_0_propagate;
    end
    if (mesh_1_1_io_out_valid_0) begin
      _T_266 <= mesh_1_1_io_out_control_0_shift;
    end
    if (mesh_1_1_io_out_valid_0) begin
      _T_268 <= mesh_1_1_io_out_control_0_propagate;
    end
    if (mesh_2_1_io_out_valid_0) begin
      _T_269 <= mesh_2_1_io_out_control_0_shift;
    end
    if (mesh_2_1_io_out_valid_0) begin
      _T_271 <= mesh_2_1_io_out_control_0_propagate;
    end
    if (mesh_3_1_io_out_valid_0) begin
      _T_272 <= mesh_3_1_io_out_control_0_shift;
    end
    if (mesh_3_1_io_out_valid_0) begin
      _T_274 <= mesh_3_1_io_out_control_0_propagate;
    end
    if (mesh_4_1_io_out_valid_0) begin
      _T_275 <= mesh_4_1_io_out_control_0_shift;
    end
    if (mesh_4_1_io_out_valid_0) begin
      _T_277 <= mesh_4_1_io_out_control_0_propagate;
    end
    if (mesh_5_1_io_out_valid_0) begin
      _T_278 <= mesh_5_1_io_out_control_0_shift;
    end
    if (mesh_5_1_io_out_valid_0) begin
      _T_280 <= mesh_5_1_io_out_control_0_propagate;
    end
    if (mesh_6_1_io_out_valid_0) begin
      _T_281 <= mesh_6_1_io_out_control_0_shift;
    end
    if (mesh_6_1_io_out_valid_0) begin
      _T_283 <= mesh_6_1_io_out_control_0_propagate;
    end
    //_T_284_0_propagate <= io_in_control_2_0_propagate;
    //_T_284_0_shift <= io_in_control_2_0_shift;
    //_T_285_0 <= io_in_valid_2_0;
     if (io_in_valid_2_0) begin
    _T_286 <= io_in_control_2_0_shift;
    end
     if (io_in_valid_2_0) begin
    _T_288 <= io_in_control_2_0_propagate;
    end
    if (mesh_0_2_io_out_valid_0) begin
      _T_289 <= mesh_0_2_io_out_control_0_shift;
    end
    if (mesh_0_2_io_out_valid_0) begin
      _T_291 <= mesh_0_2_io_out_control_0_propagate;
    end
    if (mesh_1_2_io_out_valid_0) begin
      _T_292 <= mesh_1_2_io_out_control_0_shift;
    end
    if (mesh_1_2_io_out_valid_0) begin
      _T_294 <= mesh_1_2_io_out_control_0_propagate;
    end
    if (mesh_2_2_io_out_valid_0) begin
      _T_295 <= mesh_2_2_io_out_control_0_shift;
    end
    if (mesh_2_2_io_out_valid_0) begin
      _T_297 <= mesh_2_2_io_out_control_0_propagate;
    end
    if (mesh_3_2_io_out_valid_0) begin
      _T_298 <= mesh_3_2_io_out_control_0_shift;
    end
    if (mesh_3_2_io_out_valid_0) begin
      _T_300 <= mesh_3_2_io_out_control_0_propagate;
    end
    if (mesh_4_2_io_out_valid_0) begin
      _T_301 <= mesh_4_2_io_out_control_0_shift;
    end
    if (mesh_4_2_io_out_valid_0) begin
      _T_303 <= mesh_4_2_io_out_control_0_propagate;
    end
    if (mesh_5_2_io_out_valid_0) begin
      _T_304 <= mesh_5_2_io_out_control_0_shift;
    end
    if (mesh_5_2_io_out_valid_0) begin
      _T_306 <= mesh_5_2_io_out_control_0_propagate;
    end
    if (mesh_6_2_io_out_valid_0) begin
      _T_307 <= mesh_6_2_io_out_control_0_shift;
    end
    if (mesh_6_2_io_out_valid_0) begin
      _T_309 <= mesh_6_2_io_out_control_0_propagate;
    end
    //_T_310_0_propagate <= io_in_control_3_0_propagate;
    //_T_310_0_shift <= io_in_control_3_0_shift;
    //_T_311_0 <= io_in_valid_3_0;
     if (io_in_valid_3_0) begin
    _T_312 <= io_in_control_3_0_shift;
    end
     if (io_in_valid_3_0) begin
    _T_314 <= io_in_control_3_0_propagate;
    end
    if (mesh_0_3_io_out_valid_0) begin
      _T_315 <= mesh_0_3_io_out_control_0_shift;
    end
    if (mesh_0_3_io_out_valid_0) begin
      _T_317 <= mesh_0_3_io_out_control_0_propagate;
    end
    if (mesh_1_3_io_out_valid_0) begin
      _T_318 <= mesh_1_3_io_out_control_0_shift;
    end
    if (mesh_1_3_io_out_valid_0) begin
      _T_320 <= mesh_1_3_io_out_control_0_propagate;
    end
    if (mesh_2_3_io_out_valid_0) begin
      _T_321 <= mesh_2_3_io_out_control_0_shift;
    end
    if (mesh_2_3_io_out_valid_0) begin
      _T_323 <= mesh_2_3_io_out_control_0_propagate;
    end
    if (mesh_3_3_io_out_valid_0) begin
      _T_324 <= mesh_3_3_io_out_control_0_shift;
    end
    if (mesh_3_3_io_out_valid_0) begin
      _T_326 <= mesh_3_3_io_out_control_0_propagate;
    end
    if (mesh_4_3_io_out_valid_0) begin
      _T_327 <= mesh_4_3_io_out_control_0_shift;
    end
    if (mesh_4_3_io_out_valid_0) begin
      _T_329 <= mesh_4_3_io_out_control_0_propagate;
    end
    if (mesh_5_3_io_out_valid_0) begin
      _T_330 <= mesh_5_3_io_out_control_0_shift;
    end
    if (mesh_5_3_io_out_valid_0) begin
      _T_332 <= mesh_5_3_io_out_control_0_propagate;
    end
    if (mesh_6_3_io_out_valid_0) begin
      _T_333 <= mesh_6_3_io_out_control_0_shift;
    end
    if (mesh_6_3_io_out_valid_0) begin
      _T_335 <= mesh_6_3_io_out_control_0_propagate;
    end
    //_T_336_0_propagate <= io_in_control_4_0_propagate;
    //_T_336_0_shift <= io_in_control_4_0_shift;
    //_T_337_0 <= io_in_valid_4_0;
     if (io_in_valid_4_0) begin
    _T_338 <= io_in_control_4_0_shift;
    end
     if (io_in_valid_4_0) begin
    _T_340 <= io_in_control_4_0_propagate;
    end
    if (mesh_0_4_io_out_valid_0) begin
      _T_341 <= mesh_0_4_io_out_control_0_shift;
    end
    if (mesh_0_4_io_out_valid_0) begin
      _T_343 <= mesh_0_4_io_out_control_0_propagate;
    end
    if (mesh_1_4_io_out_valid_0) begin
      _T_344 <= mesh_1_4_io_out_control_0_shift;
    end
    if (mesh_1_4_io_out_valid_0) begin
      _T_346 <= mesh_1_4_io_out_control_0_propagate;
    end
    if (mesh_2_4_io_out_valid_0) begin
      _T_347 <= mesh_2_4_io_out_control_0_shift;
    end
    if (mesh_2_4_io_out_valid_0) begin
      _T_349 <= mesh_2_4_io_out_control_0_propagate;
    end
    if (mesh_3_4_io_out_valid_0) begin
      _T_350 <= mesh_3_4_io_out_control_0_shift;
    end
    if (mesh_3_4_io_out_valid_0) begin
      _T_352 <= mesh_3_4_io_out_control_0_propagate;
    end
    if (mesh_4_4_io_out_valid_0) begin
      _T_353 <= mesh_4_4_io_out_control_0_shift;
    end
    if (mesh_4_4_io_out_valid_0) begin
      _T_355 <= mesh_4_4_io_out_control_0_propagate;
    end
    if (mesh_5_4_io_out_valid_0) begin
      _T_356 <= mesh_5_4_io_out_control_0_shift;
    end
    if (mesh_5_4_io_out_valid_0) begin
      _T_358 <= mesh_5_4_io_out_control_0_propagate;
    end
    if (mesh_6_4_io_out_valid_0) begin
      _T_359 <= mesh_6_4_io_out_control_0_shift;
    end
    if (mesh_6_4_io_out_valid_0) begin
      _T_361 <= mesh_6_4_io_out_control_0_propagate;
    end
    //_T_362_0_propagate <= io_in_control_5_0_propagate;
    //_T_362_0_shift <= io_in_control_5_0_shift;
    //_T_363_0 <= io_in_valid_5_0;
     if (io_in_valid_5_0) begin
    _T_364 <= io_in_control_5_0_shift;
    end
     if (io_in_valid_5_0) begin
    _T_366 <= io_in_control_5_0_propagate;
    end
    if (mesh_0_5_io_out_valid_0) begin
      _T_367 <= mesh_0_5_io_out_control_0_shift;
    end
    if (mesh_0_5_io_out_valid_0) begin
      _T_369 <= mesh_0_5_io_out_control_0_propagate;
    end
    if (mesh_1_5_io_out_valid_0) begin
      _T_370 <= mesh_1_5_io_out_control_0_shift;
    end
    if (mesh_1_5_io_out_valid_0) begin
      _T_372 <= mesh_1_5_io_out_control_0_propagate;
    end
    if (mesh_2_5_io_out_valid_0) begin
      _T_373 <= mesh_2_5_io_out_control_0_shift;
    end
    if (mesh_2_5_io_out_valid_0) begin
      _T_375 <= mesh_2_5_io_out_control_0_propagate;
    end
    if (mesh_3_5_io_out_valid_0) begin
      _T_376 <= mesh_3_5_io_out_control_0_shift;
    end
    if (mesh_3_5_io_out_valid_0) begin
      _T_378 <= mesh_3_5_io_out_control_0_propagate;
    end
    if (mesh_4_5_io_out_valid_0) begin
      _T_379 <= mesh_4_5_io_out_control_0_shift;
    end
    if (mesh_4_5_io_out_valid_0) begin
      _T_381 <= mesh_4_5_io_out_control_0_propagate;
    end
    if (mesh_5_5_io_out_valid_0) begin
      _T_382 <= mesh_5_5_io_out_control_0_shift;
    end
    if (mesh_5_5_io_out_valid_0) begin
      _T_384 <= mesh_5_5_io_out_control_0_propagate;
    end
    if (mesh_6_5_io_out_valid_0) begin
      _T_385 <= mesh_6_5_io_out_control_0_shift;
    end
    if (mesh_6_5_io_out_valid_0) begin
      _T_387 <= mesh_6_5_io_out_control_0_propagate;
    end
    //_T_388_0_propagate <= io_in_control_6_0_propagate;
    //_T_388_0_shift <= io_in_control_6_0_shift;
    //_T_389_0 <= io_in_valid_6_0;
     if (io_in_valid_6_0) begin
    _T_390 <= io_in_control_6_0_shift;
    end
     if (io_in_valid_6_0) begin
    _T_392 <= io_in_control_6_0_propagate;
    end
    if (mesh_0_6_io_out_valid_0) begin
      _T_393 <= mesh_0_6_io_out_control_0_shift;
    end
    if (mesh_0_6_io_out_valid_0) begin
      _T_395 <= mesh_0_6_io_out_control_0_propagate;
    end
    if (mesh_1_6_io_out_valid_0) begin
      _T_396 <= mesh_1_6_io_out_control_0_shift;
    end
    if (mesh_1_6_io_out_valid_0) begin
      _T_398 <= mesh_1_6_io_out_control_0_propagate;
    end
    if (mesh_2_6_io_out_valid_0) begin
      _T_399 <= mesh_2_6_io_out_control_0_shift;
    end
    if (mesh_2_6_io_out_valid_0) begin
      _T_401 <= mesh_2_6_io_out_control_0_propagate;
    end
    if (mesh_3_6_io_out_valid_0) begin
      _T_402 <= mesh_3_6_io_out_control_0_shift;
    end
    if (mesh_3_6_io_out_valid_0) begin
      _T_404 <= mesh_3_6_io_out_control_0_propagate;
    end
    if (mesh_4_6_io_out_valid_0) begin
      _T_405 <= mesh_4_6_io_out_control_0_shift;
    end
    if (mesh_4_6_io_out_valid_0) begin
      _T_407 <= mesh_4_6_io_out_control_0_propagate;
    end
    if (mesh_5_6_io_out_valid_0) begin
      _T_408 <= mesh_5_6_io_out_control_0_shift;
    end
    if (mesh_5_6_io_out_valid_0) begin
      _T_410 <= mesh_5_6_io_out_control_0_propagate;
    end
    if (mesh_6_6_io_out_valid_0) begin
      _T_411 <= mesh_6_6_io_out_control_0_shift;
    end
    if (mesh_6_6_io_out_valid_0) begin
      _T_413 <= mesh_6_6_io_out_control_0_propagate;
    end
    //_T_414_0_propagate <= io_in_control_7_0_propagate;
    //_T_414_0_shift <= io_in_control_7_0_shift;
    //_T_415_0 <= io_in_valid_7_0;
     if (io_in_valid_7_0) begin
    _T_416 <= io_in_control_7_0_shift;
    end
     if (io_in_valid_7_0) begin
    _T_418 <= io_in_control_7_0_propagate;
    end
    if (mesh_0_7_io_out_valid_0) begin
      _T_419 <= mesh_0_7_io_out_control_0_shift;
    end
    if (mesh_0_7_io_out_valid_0) begin
      _T_421 <= mesh_0_7_io_out_control_0_propagate;
    end
    if (mesh_1_7_io_out_valid_0) begin
      _T_422 <= mesh_1_7_io_out_control_0_shift;
    end
    if (mesh_1_7_io_out_valid_0) begin
      _T_424 <= mesh_1_7_io_out_control_0_propagate;
    end
    if (mesh_2_7_io_out_valid_0) begin
      _T_425 <= mesh_2_7_io_out_control_0_shift;
    end
    if (mesh_2_7_io_out_valid_0) begin
      _T_427 <= mesh_2_7_io_out_control_0_propagate;
    end
    if (mesh_3_7_io_out_valid_0) begin
      _T_428 <= mesh_3_7_io_out_control_0_shift;
    end
    if (mesh_3_7_io_out_valid_0) begin
      _T_430 <= mesh_3_7_io_out_control_0_propagate;
    end
    if (mesh_4_7_io_out_valid_0) begin
      _T_431 <= mesh_4_7_io_out_control_0_shift;
    end
    if (mesh_4_7_io_out_valid_0) begin
      _T_433 <= mesh_4_7_io_out_control_0_propagate;
    end
    if (mesh_5_7_io_out_valid_0) begin
      _T_434 <= mesh_5_7_io_out_control_0_shift;
    end
    if (mesh_5_7_io_out_valid_0) begin
      _T_436 <= mesh_5_7_io_out_control_0_propagate;
    end
    if (mesh_6_7_io_out_valid_0) begin
      _T_437 <= mesh_6_7_io_out_control_0_shift;
    end
    if (mesh_6_7_io_out_valid_0) begin
      _T_439 <= mesh_6_7_io_out_control_0_propagate;
    end
    //_T_440_0 <= io_in_valid_0_0;
    _T_441_0 <= io_in_valid_0_0;
    _T_442_0 <= mesh_0_0_io_out_valid_0;
    _T_443_0 <= mesh_1_0_io_out_valid_0;
    _T_444_0 <= mesh_2_0_io_out_valid_0;
    _T_445_0 <= mesh_3_0_io_out_valid_0;
    _T_446_0 <= mesh_4_0_io_out_valid_0;
    _T_447_0 <= mesh_5_0_io_out_valid_0;
    _T_448_0 <= mesh_6_0_io_out_valid_0;
    //_T_449_0 <= io_in_valid_1_0;
    _T_450_0 <= io_in_valid_1_0;
    _T_451_0 <= mesh_0_1_io_out_valid_0;
    _T_452_0 <= mesh_1_1_io_out_valid_0;
    _T_453_0 <= mesh_2_1_io_out_valid_0;
    _T_454_0 <= mesh_3_1_io_out_valid_0;
    _T_455_0 <= mesh_4_1_io_out_valid_0;
    _T_456_0 <= mesh_5_1_io_out_valid_0;
    _T_457_0 <= mesh_6_1_io_out_valid_0;
    //_T_458_0 <= io_in_valid_2_0;
    _T_459_0 <= io_in_valid_2_0;
    _T_460_0 <= mesh_0_2_io_out_valid_0;
    _T_461_0 <= mesh_1_2_io_out_valid_0;
    _T_462_0 <= mesh_2_2_io_out_valid_0;
    _T_463_0 <= mesh_3_2_io_out_valid_0;
    _T_464_0 <= mesh_4_2_io_out_valid_0;
    _T_465_0 <= mesh_5_2_io_out_valid_0;
    _T_466_0 <= mesh_6_2_io_out_valid_0;
    //_T_467_0 <= io_in_valid_3_0;
    _T_468_0 <= io_in_valid_3_0;
    _T_469_0 <= mesh_0_3_io_out_valid_0;
    _T_470_0 <= mesh_1_3_io_out_valid_0;
    _T_471_0 <= mesh_2_3_io_out_valid_0;
    _T_472_0 <= mesh_3_3_io_out_valid_0;
    _T_473_0 <= mesh_4_3_io_out_valid_0;
    _T_474_0 <= mesh_5_3_io_out_valid_0;
    _T_475_0 <= mesh_6_3_io_out_valid_0;
    //_T_476_0 <= io_in_valid_4_0;
    _T_477_0 <= io_in_valid_4_0;
    _T_478_0 <= mesh_0_4_io_out_valid_0;
    _T_479_0 <= mesh_1_4_io_out_valid_0;
    _T_480_0 <= mesh_2_4_io_out_valid_0;
    _T_481_0 <= mesh_3_4_io_out_valid_0;
    _T_482_0 <= mesh_4_4_io_out_valid_0;
    _T_483_0 <= mesh_5_4_io_out_valid_0;
    _T_484_0 <= mesh_6_4_io_out_valid_0;
    //_T_485_0 <= io_in_valid_5_0;
    _T_486_0 <= io_in_valid_5_0;
    _T_487_0 <= mesh_0_5_io_out_valid_0;
    _T_488_0 <= mesh_1_5_io_out_valid_0;
    _T_489_0 <= mesh_2_5_io_out_valid_0;
    _T_490_0 <= mesh_3_5_io_out_valid_0;
    _T_491_0 <= mesh_4_5_io_out_valid_0;
    _T_492_0 <= mesh_5_5_io_out_valid_0;
    _T_493_0 <= mesh_6_5_io_out_valid_0;
    //_T_494_0 <= io_in_valid_6_0;
    _T_495_0 <= io_in_valid_6_0;
    _T_496_0 <= mesh_0_6_io_out_valid_0;
    _T_497_0 <= mesh_1_6_io_out_valid_0;
    _T_498_0 <= mesh_2_6_io_out_valid_0;
    _T_499_0 <= mesh_3_6_io_out_valid_0;
    _T_500_0 <= mesh_4_6_io_out_valid_0;
    _T_501_0 <= mesh_5_6_io_out_valid_0;
    _T_502_0 <= mesh_6_6_io_out_valid_0;
    //_T_503_0 <= io_in_valid_7_0;
    _T_504_0 <= io_in_valid_7_0;
    _T_505_0 <= mesh_0_7_io_out_valid_0;
    _T_506_0 <= mesh_1_7_io_out_valid_0;
    _T_507_0 <= mesh_2_7_io_out_valid_0;
    _T_508_0 <= mesh_3_7_io_out_valid_0;
    _T_509_0 <= mesh_4_7_io_out_valid_0;
    _T_510_0 <= mesh_5_7_io_out_valid_0;
    _T_511_0 <= mesh_6_7_io_out_valid_0;
  end
endmodule
//////////////////////////Round/Shift////////////////////////////////////////////////////////
  module rounding(
input         clock,
input [63:0] c1,
input  [5:0]  io_in_control_shift,
input io_in_control_propagate,
input         io_in_valid,
output [18:0] _T_35
 );

  wire  last_s; // @[Reg.scala 15:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166246.4]
  wire  flip; // @[PE.scala 58:21:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166250.4]
  wire [5:0] shift_offset; // @[PE.scala 59:25:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166251.4]
  wire  _T_4; // @[Arithmetic.scala 72:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166258.8]
  wire [5:0] _T_6; // @[Arithmetic.scala 72:53:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166260.8]
  wire [63:0] _T_7; // @[Arithmetic.scala 72:50:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166261.8]
  wire  _T_8; // @[Arithmetic.scala 72:50:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166262.8]
  wire  _T_9; // @[Arithmetic.scala 72:29:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166263.8]
  wire  _T_10; // @[Arithmetic.scala 73:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166264.8]
  wire [63:0] _T_11; // @[Arithmetic.scala 73:51:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166265.8]
  wire [63:0] _T_14; // @[Arithmetic.scala 73:62:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166268.8]
  wire [63:0] _T_16; // @[Arithmetic.scala 73:85:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166270.8]
  wire [63:0] _T_17; // @[Arithmetic.scala 73:54:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166271.8]
  wire [63:0] _T_18; // @[Arithmetic.scala 73:24:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166272.8]
  wire  _T_19; // @[Arithmetic.scala 73:93:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166273.8]
  wire [63:0] _T_20; // @[Arithmetic.scala 74:30:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166274.8]
  wire  _T_21; // @[Arithmetic.scala 74:30:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166275.8]
  wire  _T_22; // @[Arithmetic.scala 76:38:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166276.8]
  wire  _T_23; // @[Arithmetic.scala 76:29:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166277.8]
  wire [1:0] _T_26; // @[Arithmetic.scala 78:35:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166280.8]
  wire [63:0] _GEN_19; // @[Arithmetic.scala 78:30:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166281.8]
  wire [63:0] _T_28; // @[Arithmetic.scala 78:30:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166282.8]
  wire [63:0] _T_29; // @[Arithmetic.scala 78:30:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166283.8]
  wire  _T_30; // @[Arithmetic.scala 86:33:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166284.8]
  wire  _T_31; // @[Arithmetic.scala 86:60:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166285.8]
  wire [63:0] _T_32; // @[Mux.scala 87:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166286.8]
  wire [63:0] _T_33; // @[Mux.scala 87:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166287.8]
  wire [18:0] _T_34; // @[Arithmetic.scala 86:81:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166288.8]
  //wire [18:0] _T_35; // @[Arithmetic.scala 86:105:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166289.8]

  assign last_s =io_in_control_propagate;
  assign flip = last_s != io_in_control_propagate; // @[PE.scala 58:21:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166250.4]
  assign shift_offset = flip ? io_in_control_shift : 6'h0; // @[PE.scala 59:25:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166251.4]
  assign _T_4 = shift_offset == 6'h0; // @[Arithmetic.scala 72:32:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166258.8]
  assign _T_6 = shift_offset - 6'h1; // @[Arithmetic.scala 72:53:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166260.8]
  assign _T_7 = $signed(c1) >>> _T_6; // @[Arithmetic.scala 72:50:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166261.8]
  assign _T_8 = _T_7[0]; // @[Arithmetic.scala 72:50:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166262.8]
  assign _T_9 = _T_4 ? 1'h0 : _T_8; // @[Arithmetic.scala 72:29:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166263.8]
  assign _T_10 = shift_offset <= 6'h1; // @[Arithmetic.scala 73:27:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166264.8]
  assign _T_11 = $unsigned(c1); // @[Arithmetic.scala 73:51:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166265.8]
  assign _T_14 = 64'h1 << _T_6; // @[Arithmetic.scala 73:62:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166268.8]
  assign _T_16 = _T_14 - 64'h1; // @[Arithmetic.scala 73:85:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166270.8]
  assign _T_17 = _T_11 & _T_16; // @[Arithmetic.scala 73:54:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166271.8]
  assign _T_18 = _T_10 ? 64'h0 : _T_17; // @[Arithmetic.scala 73:24:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166272.8]
  assign _T_19 = _T_18 != 64'h0; // @[Arithmetic.scala 73:93:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166273.8]
  assign _T_20 = $signed(c1) >>> shift_offset; // @[Arithmetic.scala 74:30:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166274.8]
  assign _T_21 = _T_20[0]; // @[Arithmetic.scala 74:30:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166275.8]
  assign _T_22 = _T_19 | _T_21; // @[Arithmetic.scala 76:38:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166276.8]
  assign _T_23 = _T_9 & _T_22; // @[Arithmetic.scala 76:29:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166277.8]
  assign _T_26 = _T_23 ? $signed(2'sh1) : $signed(2'sh0); // @[Arithmetic.scala 78:35:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166280.8]
  assign _GEN_19 = {{62{_T_26[1]}},_T_26}; // @[Arithmetic.scala 78:30:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166281.8]
  assign _T_28 = $signed(_T_20) + $signed(_GEN_19); // @[Arithmetic.scala 78:30:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166282.8]
  assign _T_29 = $signed(_T_28); // @[Arithmetic.scala 78:30:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166283.8]
  assign _T_30 = $signed(_T_29) > $signed(64'sh3ffff); // @[Arithmetic.scala 86:33:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166284.8]
  assign _T_31 = $signed(_T_29) < $signed(-64'sh40000); // @[Arithmetic.scala 86:60:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166285.8]
  assign _T_32 = _T_31 ? $signed(-64'sh40000) : $signed(_T_29); // @[Mux.scala 87:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166286.8]
  assign _T_33 = _T_30 ? $signed(64'sh3ffff) : $signed(_T_32); // @[Mux.scala 87:16:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166287.8]
  assign _T_34 = _T_33[18:0]; // @[Arithmetic.scala 86:81:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166288.8]
  assign _T_35 = $signed(_T_34); // @[Arithmetic.scala 86:105:example.TestHarness.GemminiSocTest1RocketConfig864.fir@166289.8]
  endmodule